magic
tech sky130A
magscale 1 2
timestamp 1608250781
<< viali >>
rect 4813 12257 4847 12291
rect 8217 12257 8251 12291
rect 4537 12189 4571 12223
rect 5917 12053 5951 12087
rect 8309 12053 8343 12087
rect 2697 11713 2731 11747
rect 4721 11713 4755 11747
rect 7573 11713 7607 11747
rect 2973 11645 3007 11679
rect 4445 11645 4479 11679
rect 7665 11645 7699 11679
rect 8125 11577 8159 11611
rect 4261 11509 4295 11543
rect 6009 11509 6043 11543
rect 10701 11305 10735 11339
rect 4077 11169 4111 11203
rect 4353 11169 4387 11203
rect 6285 11169 6319 11203
rect 7665 11169 7699 11203
rect 7757 11169 7791 11203
rect 10609 11169 10643 11203
rect 5549 11101 5583 11135
rect 6837 11101 6871 11135
rect 6929 11101 6963 11135
rect 6377 10965 6411 10999
rect 7803 10761 7837 10795
rect 8309 10761 8343 10795
rect 7941 10693 7975 10727
rect 5365 10625 5399 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 8033 10625 8067 10659
rect 5917 10557 5951 10591
rect 6193 10557 6227 10591
rect 6469 10557 6503 10591
rect 6837 10557 6871 10591
rect 7297 10557 7331 10591
rect 7573 10557 7607 10591
rect 7665 10489 7699 10523
rect 4629 10217 4663 10251
rect 2973 10149 3007 10183
rect 8769 10149 8803 10183
rect 2513 10081 2547 10115
rect 4537 10081 4571 10115
rect 4813 10081 4847 10115
rect 4905 10081 4939 10115
rect 5089 10081 5123 10115
rect 5733 10081 5767 10115
rect 6193 10081 6227 10115
rect 6561 10081 6595 10115
rect 7389 10081 7423 10115
rect 7665 10081 7699 10115
rect 7941 10081 7975 10115
rect 8953 10081 8987 10115
rect 2421 10013 2455 10047
rect 5273 10013 5307 10047
rect 6837 10013 6871 10047
rect 7849 10013 7883 10047
rect 8309 10013 8343 10047
rect 6469 9945 6503 9979
rect 8106 9945 8140 9979
rect 8217 9877 8251 9911
rect 8585 9877 8619 9911
rect 9045 9877 9079 9911
rect 7113 9673 7147 9707
rect 4445 9605 4479 9639
rect 3893 9537 3927 9571
rect 6285 9537 6319 9571
rect 7757 9537 7791 9571
rect 8125 9537 8159 9571
rect 9137 9537 9171 9571
rect 9965 9537 9999 9571
rect 1409 9469 1443 9503
rect 3801 9469 3835 9503
rect 4077 9469 4111 9503
rect 4629 9469 4663 9503
rect 5089 9469 5123 9503
rect 5641 9469 5675 9503
rect 5825 9469 5859 9503
rect 6009 9469 6043 9503
rect 6653 9469 6687 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 7849 9469 7883 9503
rect 8677 9469 8711 9503
rect 8953 9469 8987 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 9873 9469 9907 9503
rect 5181 9401 5215 9435
rect 9781 9401 9815 9435
rect 1501 9333 1535 9367
rect 4169 9333 4203 9367
rect 2329 9129 2363 9163
rect 3525 9129 3559 9163
rect 9781 9129 9815 9163
rect 10609 9129 10643 9163
rect 5089 9061 5123 9095
rect 1869 8993 1903 9027
rect 2237 8993 2271 9027
rect 3433 8993 3467 9027
rect 3709 8993 3743 9027
rect 4261 8993 4295 9027
rect 4997 8993 5031 9027
rect 5549 8993 5583 9027
rect 5733 8993 5767 9027
rect 6101 8993 6135 9027
rect 6837 8993 6871 9027
rect 7021 8993 7055 9027
rect 7205 8993 7239 9027
rect 7941 8993 7975 9027
rect 8769 8993 8803 9027
rect 9045 8993 9079 9027
rect 9689 8993 9723 9027
rect 10149 8993 10183 9027
rect 10517 8993 10551 9027
rect 10793 8993 10827 9027
rect 6009 8925 6043 8959
rect 6377 8925 6411 8959
rect 7665 8925 7699 8959
rect 7757 8925 7791 8959
rect 8493 8925 8527 8959
rect 8953 8925 8987 8959
rect 2053 8789 2087 8823
rect 3801 8789 3835 8823
rect 4353 8789 4387 8823
rect 9229 8789 9263 8823
rect 10885 8789 10919 8823
rect 3433 8585 3467 8619
rect 10885 8585 10919 8619
rect 4445 8449 4479 8483
rect 5457 8449 5491 8483
rect 7941 8449 7975 8483
rect 8217 8449 8251 8483
rect 2145 8381 2179 8415
rect 2329 8381 2363 8415
rect 2651 8381 2685 8415
rect 2789 8381 2823 8415
rect 3341 8381 3375 8415
rect 3617 8381 3651 8415
rect 3709 8381 3743 8415
rect 3893 8381 3927 8415
rect 4353 8381 4387 8415
rect 4997 8381 5031 8415
rect 5273 8381 5307 8415
rect 5549 8381 5583 8415
rect 5917 8381 5951 8415
rect 6377 8381 6411 8415
rect 6653 8381 6687 8415
rect 7297 8381 7331 8415
rect 7481 8381 7515 8415
rect 7665 8381 7699 8415
rect 8953 8381 8987 8415
rect 9229 8381 9263 8415
rect 9413 8381 9447 8415
rect 10057 8381 10091 8415
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 6837 8313 6871 8347
rect 8401 8313 8435 8347
rect 9505 8313 9539 8347
rect 1961 8245 1995 8279
rect 2789 8041 2823 8075
rect 10977 8041 11011 8075
rect 2145 7973 2179 8007
rect 5365 7973 5399 8007
rect 2292 7905 2326 7939
rect 4353 7905 4387 7939
rect 4813 7905 4847 7939
rect 5089 7905 5123 7939
rect 5825 7905 5859 7939
rect 6101 7905 6135 7939
rect 6285 7905 6319 7939
rect 7481 7905 7515 7939
rect 7573 7905 7607 7939
rect 7849 7905 7883 7939
rect 8585 7905 8619 7939
rect 9689 7905 9723 7939
rect 9919 7905 9953 7939
rect 10517 7905 10551 7939
rect 10793 7905 10827 7939
rect 2513 7837 2547 7871
rect 4445 7837 4479 7871
rect 5273 7837 5307 7871
rect 6469 7837 6503 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 8861 7837 8895 7871
rect 10057 7837 10091 7871
rect 10149 7769 10183 7803
rect 2421 7701 2455 7735
rect 9827 7701 9861 7735
rect 10609 7701 10643 7735
rect 6929 7497 6963 7531
rect 8861 7429 8895 7463
rect 4353 7361 4387 7395
rect 5365 7361 5399 7395
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 4997 7293 5031 7327
rect 5917 7293 5951 7327
rect 6101 7293 6135 7327
rect 6469 7293 6503 7327
rect 6561 7293 6595 7327
rect 6837 7293 6871 7327
rect 7757 7293 7791 7327
rect 7941 7293 7975 7327
rect 8125 7293 8159 7327
rect 8493 7293 8527 7327
rect 8677 7293 8711 7327
rect 8861 7293 8895 7327
rect 9321 7293 9355 7327
rect 9597 7293 9631 7327
rect 9873 7293 9907 7327
rect 4629 7225 4663 7259
rect 4813 7225 4847 7259
rect 7205 7225 7239 7259
rect 5733 7157 5767 7191
rect 9689 7157 9723 7191
rect 9965 7157 9999 7191
rect 9045 6953 9079 6987
rect 5457 6885 5491 6919
rect 4905 6817 4939 6851
rect 4997 6817 5031 6851
rect 6193 6817 6227 6851
rect 6561 6817 6595 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 8401 6817 8435 6851
rect 8769 6817 8803 6851
rect 8953 6817 8987 6851
rect 9873 6817 9907 6851
rect 6009 6749 6043 6783
rect 6469 6749 6503 6783
rect 6837 6749 6871 6783
rect 7389 6749 7423 6783
rect 7849 6749 7883 6783
rect 8585 6749 8619 6783
rect 5825 6613 5859 6647
rect 9965 6613 9999 6647
rect 5917 6409 5951 6443
rect 7941 6409 7975 6443
rect 10701 6409 10735 6443
rect 6561 6273 6595 6307
rect 8401 6273 8435 6307
rect 5641 6205 5675 6239
rect 6101 6205 6135 6239
rect 6285 6205 6319 6239
rect 6837 6205 6871 6239
rect 6929 6205 6963 6239
rect 7113 6205 7147 6239
rect 7665 6205 7699 6239
rect 7849 6205 7883 6239
rect 8309 6205 8343 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 9689 6205 9723 6239
rect 9873 6205 9907 6239
rect 10425 6205 10459 6239
rect 10609 6205 10643 6239
rect 7573 6137 7607 6171
rect 10149 6069 10183 6103
rect 6377 5865 6411 5899
rect 7665 5865 7699 5899
rect 7481 5797 7515 5831
rect 7941 5797 7975 5831
rect 6285 5729 6319 5763
rect 6745 5729 6779 5763
rect 7205 5729 7239 5763
rect 7573 5729 7607 5763
rect 7849 5729 7883 5763
rect 10333 5729 10367 5763
rect 10701 5729 10735 5763
rect 9689 5661 9723 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 1409 4641 1443 4675
rect 1593 4437 1627 4471
rect 10885 3689 10919 3723
rect 9873 3553 9907 3587
rect 10333 3553 10367 3587
rect 10425 3553 10459 3587
rect 9781 3485 9815 3519
rect 10241 3145 10275 3179
rect 9137 3077 9171 3111
rect 9321 2941 9355 2975
rect 9505 2941 9539 2975
rect 9873 2941 9907 2975
rect 9965 2941 9999 2975
rect 10149 2941 10183 2975
rect 10057 2601 10091 2635
rect 8217 2465 8251 2499
rect 8585 2465 8619 2499
rect 9781 2465 9815 2499
rect 9965 2465 9999 2499
rect 8309 2261 8343 2295
rect 8769 2261 8803 2295
<< metal1 >>
rect 1104 12538 11684 12560
rect 1104 12486 4508 12538
rect 4560 12486 4572 12538
rect 4624 12486 4636 12538
rect 4688 12486 4700 12538
rect 4752 12486 8035 12538
rect 8087 12486 8099 12538
rect 8151 12486 8163 12538
rect 8215 12486 8227 12538
rect 8279 12486 11684 12538
rect 1104 12464 11684 12486
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5718 12288 5724 12300
rect 4847 12260 5724 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8938 12288 8944 12300
rect 8251 12260 8944 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4120 12192 4537 12220
rect 4120 12180 4126 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 5905 12087 5963 12093
rect 5905 12084 5917 12087
rect 5500 12056 5917 12084
rect 5500 12044 5506 12056
rect 5905 12053 5917 12056
rect 5951 12053 5963 12087
rect 5905 12047 5963 12053
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 7708 12056 8309 12084
rect 7708 12044 7714 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 8297 12047 8355 12053
rect 1104 11994 11684 12016
rect 1104 11942 2745 11994
rect 2797 11942 2809 11994
rect 2861 11942 2873 11994
rect 2925 11942 2937 11994
rect 2989 11942 6272 11994
rect 6324 11942 6336 11994
rect 6388 11942 6400 11994
rect 6452 11942 6464 11994
rect 6516 11942 9798 11994
rect 9850 11942 9862 11994
rect 9914 11942 9926 11994
rect 9978 11942 9990 11994
rect 10042 11942 11684 11994
rect 1104 11920 11684 11942
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1854 11744 1860 11756
rect 1544 11716 1860 11744
rect 1544 11704 1550 11716
rect 1854 11704 1860 11716
rect 1912 11744 1918 11756
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 1912 11716 2697 11744
rect 1912 11704 1918 11716
rect 2685 11713 2697 11716
rect 2731 11744 2743 11747
rect 2731 11716 3556 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2961 11679 3019 11685
rect 2961 11676 2973 11679
rect 2832 11648 2973 11676
rect 2832 11636 2838 11648
rect 2961 11645 2973 11648
rect 3007 11645 3019 11679
rect 3528 11676 3556 11716
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 3660 11716 4721 11744
rect 3660 11704 3666 11716
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11744 7619 11747
rect 7926 11744 7932 11756
rect 7607 11716 7932 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 4062 11676 4068 11688
rect 3528 11648 4068 11676
rect 2961 11639 3019 11645
rect 4062 11636 4068 11648
rect 4120 11676 4126 11688
rect 4433 11679 4491 11685
rect 4433 11676 4445 11679
rect 4120 11648 4445 11676
rect 4120 11636 4126 11648
rect 4433 11645 4445 11648
rect 4479 11645 4491 11679
rect 7650 11676 7656 11688
rect 7611 11648 7656 11676
rect 4433 11639 4491 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8113 11611 8171 11617
rect 8113 11608 8125 11611
rect 7984 11580 8125 11608
rect 7984 11568 7990 11580
rect 8113 11577 8125 11580
rect 8159 11577 8171 11611
rect 8113 11571 8171 11577
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 5718 11540 5724 11552
rect 4295 11512 5724 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 5994 11540 6000 11552
rect 5955 11512 6000 11540
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 1104 11450 11684 11472
rect 1104 11398 4508 11450
rect 4560 11398 4572 11450
rect 4624 11398 4636 11450
rect 4688 11398 4700 11450
rect 4752 11398 8035 11450
rect 8087 11398 8099 11450
rect 8151 11398 8163 11450
rect 8215 11398 8227 11450
rect 8279 11398 11684 11450
rect 1104 11376 11684 11398
rect 10686 11336 10692 11348
rect 10647 11308 10692 11336
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7064 11240 7788 11268
rect 7064 11228 7070 11240
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4798 11200 4804 11212
rect 4387 11172 4804 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6273 11203 6331 11209
rect 6273 11200 6285 11203
rect 6144 11172 6285 11200
rect 6144 11160 6150 11172
rect 6273 11169 6285 11172
rect 6319 11169 6331 11203
rect 7650 11200 7656 11212
rect 7611 11172 7656 11200
rect 6273 11163 6331 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 7760 11209 7788 11240
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10468 11172 10609 11200
rect 10468 11160 10474 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 5534 11132 5540 11144
rect 5495 11104 5540 11132
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 8386 11132 8392 11144
rect 6963 11104 8392 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 474 11024 480 11076
rect 532 11064 538 11076
rect 1486 11064 1492 11076
rect 532 11036 1492 11064
rect 532 11024 538 11036
rect 1486 11024 1492 11036
rect 1544 11024 1550 11076
rect 6840 11064 6868 11095
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 8294 11064 8300 11076
rect 6840 11036 8300 11064
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 6365 10999 6423 11005
rect 6365 10965 6377 10999
rect 6411 10996 6423 10999
rect 6822 10996 6828 11008
rect 6411 10968 6828 10996
rect 6411 10965 6423 10968
rect 6365 10959 6423 10965
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 1104 10906 11684 10928
rect 1104 10854 2745 10906
rect 2797 10854 2809 10906
rect 2861 10854 2873 10906
rect 2925 10854 2937 10906
rect 2989 10854 6272 10906
rect 6324 10854 6336 10906
rect 6388 10854 6400 10906
rect 6452 10854 6464 10906
rect 6516 10854 9798 10906
rect 9850 10854 9862 10906
rect 9914 10854 9926 10906
rect 9978 10854 9990 10906
rect 10042 10854 11684 10906
rect 1104 10832 11684 10854
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7791 10795 7849 10801
rect 7791 10792 7803 10795
rect 7708 10764 7803 10792
rect 7708 10752 7714 10764
rect 7791 10761 7803 10764
rect 7837 10761 7849 10795
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 7791 10755 7849 10761
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 5994 10684 6000 10736
rect 6052 10724 6058 10736
rect 7929 10727 7987 10733
rect 6052 10696 6500 10724
rect 6052 10684 6058 10696
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5626 10656 5632 10668
rect 5399 10628 5632 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5626 10616 5632 10628
rect 5684 10656 5690 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5684 10628 6377 10656
rect 5684 10616 5690 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6472 10597 6500 10696
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8846 10724 8852 10736
rect 7975 10696 8852 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8846 10684 8852 10696
rect 8904 10724 8910 10736
rect 9674 10724 9680 10736
rect 8904 10696 9680 10724
rect 8904 10684 8910 10696
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 7742 10656 7748 10668
rect 6595 10628 7748 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7892 10628 8033 10656
rect 7892 10616 7898 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 5905 10591 5963 10597
rect 5905 10588 5917 10591
rect 5868 10560 5917 10588
rect 5868 10548 5874 10560
rect 5905 10557 5917 10560
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10557 6239 10591
rect 6181 10551 6239 10557
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10588 6515 10591
rect 6638 10588 6644 10600
rect 6503 10560 6644 10588
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 4890 10480 4896 10532
rect 4948 10520 4954 10532
rect 6196 10520 6224 10551
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7282 10588 7288 10600
rect 7243 10560 7288 10588
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 8754 10588 8760 10600
rect 7607 10560 8760 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 4948 10492 6224 10520
rect 4948 10480 4954 10492
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7653 10523 7711 10529
rect 7653 10520 7665 10523
rect 6972 10492 7665 10520
rect 6972 10480 6978 10492
rect 7653 10489 7665 10492
rect 7699 10489 7711 10523
rect 7653 10483 7711 10489
rect 8386 10480 8392 10532
rect 8444 10520 8450 10532
rect 9030 10520 9036 10532
rect 8444 10492 9036 10520
rect 8444 10480 8450 10492
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 9674 10452 9680 10464
rect 6880 10424 9680 10452
rect 6880 10412 6886 10424
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 1104 10362 11684 10384
rect 1104 10310 4508 10362
rect 4560 10310 4572 10362
rect 4624 10310 4636 10362
rect 4688 10310 4700 10362
rect 4752 10310 8035 10362
rect 8087 10310 8099 10362
rect 8151 10310 8163 10362
rect 8215 10310 8227 10362
rect 8279 10310 11684 10362
rect 1104 10288 11684 10310
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5074 10248 5080 10260
rect 4663 10220 5080 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5074 10208 5080 10220
rect 5132 10248 5138 10260
rect 5810 10248 5816 10260
rect 5132 10220 5816 10248
rect 5132 10208 5138 10220
rect 5810 10208 5816 10220
rect 5868 10248 5874 10260
rect 8662 10248 8668 10260
rect 5868 10220 8668 10248
rect 5868 10208 5874 10220
rect 2961 10183 3019 10189
rect 2961 10149 2973 10183
rect 3007 10180 3019 10183
rect 4062 10180 4068 10192
rect 3007 10152 4068 10180
rect 3007 10149 3019 10152
rect 2961 10143 3019 10149
rect 4062 10140 4068 10152
rect 4120 10180 4126 10192
rect 4120 10152 4936 10180
rect 4120 10140 4126 10152
rect 4908 10124 4936 10152
rect 5626 10140 5632 10192
rect 5684 10180 5690 10192
rect 5684 10152 5764 10180
rect 5684 10140 5690 10152
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4396 10084 4537 10112
rect 4396 10072 4402 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4798 10112 4804 10124
rect 4759 10084 4804 10112
rect 4525 10075 4583 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 4890 10072 4896 10124
rect 4948 10112 4954 10124
rect 5736 10121 5764 10152
rect 5077 10115 5135 10121
rect 4948 10084 4993 10112
rect 4948 10072 4954 10084
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5721 10115 5779 10121
rect 5123 10084 5672 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 3050 10044 3056 10056
rect 2455 10016 3056 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5644 9988 5672 10084
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 5810 10112 5816 10124
rect 5767 10084 5816 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10112 6607 10115
rect 6730 10112 6736 10124
rect 6595 10084 6736 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 6196 10044 6224 10075
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 7392 10121 7420 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 8757 10183 8815 10189
rect 8757 10180 8769 10183
rect 7524 10152 8769 10180
rect 7524 10140 7530 10152
rect 8757 10149 8769 10152
rect 8803 10149 8815 10183
rect 8757 10143 8815 10149
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 7650 10112 7656 10124
rect 7611 10084 7656 10112
rect 7377 10075 7435 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8386 10112 8392 10124
rect 7975 10084 8392 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8904 10084 8953 10112
rect 8904 10072 8910 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6196 10016 6837 10044
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 7006 10044 7012 10056
rect 6871 10016 7012 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7006 10004 7012 10016
rect 7064 10044 7070 10056
rect 7837 10047 7895 10053
rect 7064 10016 7604 10044
rect 7064 10004 7070 10016
rect 3418 9936 3424 9988
rect 3476 9976 3482 9988
rect 4798 9976 4804 9988
rect 3476 9948 4804 9976
rect 3476 9936 3482 9948
rect 4798 9936 4804 9948
rect 4856 9936 4862 9988
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 5684 9948 6469 9976
rect 5684 9936 5690 9948
rect 6457 9945 6469 9948
rect 6503 9945 6515 9979
rect 7576 9976 7604 10016
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 9398 10044 9404 10056
rect 8343 10016 9404 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 7852 9976 7880 10007
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 7576 9948 7880 9976
rect 8094 9979 8152 9985
rect 6457 9939 6515 9945
rect 8094 9945 8106 9979
rect 8140 9976 8152 9979
rect 8478 9976 8484 9988
rect 8140 9948 8484 9976
rect 8140 9945 8152 9948
rect 8094 9939 8152 9945
rect 8478 9936 8484 9948
rect 8536 9936 8542 9988
rect 4816 9908 4844 9936
rect 7650 9908 7656 9920
rect 4816 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 7984 9880 8217 9908
rect 7984 9868 7990 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 8938 9908 8944 9920
rect 8619 9880 8944 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 9033 9911 9091 9917
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 9122 9908 9128 9920
rect 9079 9880 9128 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 1104 9818 11684 9840
rect 1104 9766 2745 9818
rect 2797 9766 2809 9818
rect 2861 9766 2873 9818
rect 2925 9766 2937 9818
rect 2989 9766 6272 9818
rect 6324 9766 6336 9818
rect 6388 9766 6400 9818
rect 6452 9766 6464 9818
rect 6516 9766 9798 9818
rect 9850 9766 9862 9818
rect 9914 9766 9926 9818
rect 9978 9766 9990 9818
rect 10042 9766 11684 9818
rect 1104 9744 11684 9766
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 5258 9704 5264 9716
rect 3752 9676 5264 9704
rect 3752 9664 3758 9676
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 7101 9707 7159 9713
rect 7101 9704 7113 9707
rect 5500 9676 7113 9704
rect 5500 9664 5506 9676
rect 7101 9673 7113 9676
rect 7147 9704 7159 9707
rect 7282 9704 7288 9716
rect 7147 9676 7288 9704
rect 7147 9673 7159 9676
rect 7101 9667 7159 9673
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 10318 9704 10324 9716
rect 7984 9676 10324 9704
rect 7984 9664 7990 9676
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 12158 9704 12164 9716
rect 10560 9676 12164 9704
rect 10560 9664 10566 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 4433 9639 4491 9645
rect 4433 9605 4445 9639
rect 4479 9636 4491 9639
rect 10686 9636 10692 9648
rect 4479 9608 6684 9636
rect 4479 9605 4491 9608
rect 4433 9599 4491 9605
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 3927 9540 6040 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9469 3847 9503
rect 4062 9500 4068 9512
rect 4023 9472 4068 9500
rect 3789 9463 3847 9469
rect 3804 9432 3832 9463
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 4982 9500 4988 9512
rect 4663 9472 4988 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5442 9500 5448 9512
rect 5123 9472 5448 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 5810 9500 5816 9512
rect 5771 9472 5816 9500
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 6012 9509 6040 9540
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6273 9571 6331 9577
rect 6273 9568 6285 9571
rect 6144 9540 6285 9568
rect 6144 9528 6150 9540
rect 6273 9537 6285 9540
rect 6319 9537 6331 9571
rect 6273 9531 6331 9537
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 5169 9435 5227 9441
rect 3804 9404 5120 9432
rect 1489 9367 1547 9373
rect 1489 9333 1501 9367
rect 1535 9364 1547 9367
rect 2406 9364 2412 9376
rect 1535 9336 2412 9364
rect 1535 9333 1547 9336
rect 1489 9327 1547 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 4154 9364 4160 9376
rect 4115 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 5092 9364 5120 9404
rect 5169 9401 5181 9435
rect 5215 9432 5227 9435
rect 6104 9432 6132 9528
rect 6656 9509 6684 9608
rect 7760 9608 10692 9636
rect 7760 9580 7788 9608
rect 7742 9568 7748 9580
rect 7703 9540 7748 9568
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8570 9568 8576 9580
rect 8159 9540 8576 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8570 9528 8576 9540
rect 8628 9568 8634 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8628 9540 9137 9568
rect 8628 9528 8634 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 6914 9500 6920 9512
rect 6687 9472 6920 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7282 9500 7288 9512
rect 7243 9472 7288 9500
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 7484 9432 7512 9460
rect 5215 9404 6132 9432
rect 6196 9404 7512 9432
rect 7852 9432 7880 9463
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 7984 9472 8677 9500
rect 7984 9460 7990 9472
rect 8665 9469 8677 9472
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9030 9500 9036 9512
rect 8987 9472 9036 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9214 9500 9220 9512
rect 9175 9472 9220 9500
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9324 9509 9352 9608
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9548 9540 9965 9568
rect 9548 9528 9554 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10226 9500 10232 9512
rect 9907 9472 10232 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10226 9460 10232 9472
rect 10284 9500 10290 9512
rect 11054 9500 11060 9512
rect 10284 9472 11060 9500
rect 10284 9460 10290 9472
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 7852 9404 7972 9432
rect 5215 9401 5227 9404
rect 5169 9395 5227 9401
rect 5350 9364 5356 9376
rect 5092 9336 5356 9364
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 6196 9364 6224 9404
rect 5776 9336 6224 9364
rect 5776 9324 5782 9336
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 7944 9364 7972 9404
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 9769 9435 9827 9441
rect 9769 9432 9781 9435
rect 9548 9404 9781 9432
rect 9548 9392 9554 9404
rect 9769 9401 9781 9404
rect 9815 9401 9827 9435
rect 9769 9395 9827 9401
rect 10594 9364 10600 9376
rect 6328 9336 10600 9364
rect 6328 9324 6334 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 1104 9274 11684 9296
rect 1104 9222 4508 9274
rect 4560 9222 4572 9274
rect 4624 9222 4636 9274
rect 4688 9222 4700 9274
rect 4752 9222 8035 9274
rect 8087 9222 8099 9274
rect 8151 9222 8163 9274
rect 8215 9222 8227 9274
rect 8279 9222 11684 9274
rect 1104 9200 11684 9222
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2498 9160 2504 9172
rect 2363 9132 2504 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 5810 9160 5816 9172
rect 3559 9132 5816 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6822 9160 6828 9172
rect 6236 9132 6828 9160
rect 6236 9120 6242 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 9214 9160 9220 9172
rect 7340 9132 9220 9160
rect 7340 9120 7346 9132
rect 9214 9120 9220 9132
rect 9272 9160 9278 9172
rect 9490 9160 9496 9172
rect 9272 9132 9496 9160
rect 9272 9120 9278 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9129 9827 9163
rect 10594 9160 10600 9172
rect 10555 9132 10600 9160
rect 9769 9123 9827 9129
rect 5077 9095 5135 9101
rect 3436 9064 4292 9092
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 2222 9024 2228 9036
rect 2183 8996 2228 9024
rect 2222 8984 2228 8996
rect 2280 9024 2286 9036
rect 3050 9024 3056 9036
rect 2280 8996 3056 9024
rect 2280 8984 2286 8996
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3436 9033 3464 9064
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 8993 3479 9027
rect 3694 9024 3700 9036
rect 3655 8996 3700 9024
rect 3421 8987 3479 8993
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4264 9033 4292 9064
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 5166 9092 5172 9104
rect 5123 9064 5172 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5258 9052 5264 9104
rect 5316 9092 5322 9104
rect 9784 9092 9812 9123
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 10778 9120 10784 9172
rect 10836 9120 10842 9172
rect 10796 9092 10824 9120
rect 5316 9064 9812 9092
rect 9876 9064 10824 9092
rect 5316 9052 5322 9064
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4430 9024 4436 9036
rect 4295 8996 4436 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 8993 5043 9027
rect 4985 8987 5043 8993
rect 5000 8888 5028 8987
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 5500 8996 5549 9024
rect 5500 8984 5506 8996
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 6089 9027 6147 9033
rect 5767 8996 5856 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 5828 8968 5856 8996
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 6270 9024 6276 9036
rect 6135 8996 6276 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7006 9024 7012 9036
rect 6967 8996 7012 9024
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7239 8996 7941 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7929 8993 7941 8996
rect 7975 9024 7987 9027
rect 8754 9024 8760 9036
rect 7975 8996 8616 9024
rect 8715 8996 8760 9024
rect 7975 8993 7987 8996
rect 7929 8987 7987 8993
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6178 8956 6184 8968
rect 6043 8928 6184 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 6362 8956 6368 8968
rect 6323 8928 6368 8956
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7208 8956 7236 8987
rect 6788 8928 7236 8956
rect 7653 8959 7711 8965
rect 6788 8916 6794 8928
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7006 8888 7012 8900
rect 5000 8860 7012 8888
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 7668 8888 7696 8919
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8481 8959 8539 8965
rect 7800 8928 7845 8956
rect 7800 8916 7806 8928
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8588 8956 8616 8996
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9030 9024 9036 9036
rect 8991 8996 9036 9024
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 9876 9024 9904 9064
rect 9824 8996 9904 9024
rect 10137 9027 10195 9033
rect 9824 8984 9830 8996
rect 10137 8993 10149 9027
rect 10183 8993 10195 9027
rect 10502 9024 10508 9036
rect 10463 8996 10508 9024
rect 10137 8987 10195 8993
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8588 8928 8953 8956
rect 8481 8919 8539 8925
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 8202 8888 8208 8900
rect 7668 8860 8208 8888
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 8496 8888 8524 8919
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 10152 8956 10180 8987
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 9180 8928 10180 8956
rect 9180 8916 9186 8928
rect 8662 8888 8668 8900
rect 8496 8860 8668 8888
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 10796 8888 10824 8987
rect 8772 8860 10824 8888
rect 1486 8780 1492 8832
rect 1544 8820 1550 8832
rect 2041 8823 2099 8829
rect 2041 8820 2053 8823
rect 1544 8792 2053 8820
rect 1544 8780 1550 8792
rect 2041 8789 2053 8792
rect 2087 8789 2099 8823
rect 2041 8783 2099 8789
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3660 8792 3801 8820
rect 3660 8780 3666 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 7466 8820 7472 8832
rect 4387 8792 7472 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 8772 8820 8800 8860
rect 7616 8792 8800 8820
rect 7616 8780 7622 8792
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9030 8820 9036 8832
rect 8904 8792 9036 8820
rect 8904 8780 8910 8792
rect 9030 8780 9036 8792
rect 9088 8820 9094 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 9088 8792 9229 8820
rect 9088 8780 9094 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 9364 8792 10885 8820
rect 9364 8780 9370 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 10873 8783 10931 8789
rect 1104 8730 11684 8752
rect 1104 8678 2745 8730
rect 2797 8678 2809 8730
rect 2861 8678 2873 8730
rect 2925 8678 2937 8730
rect 2989 8678 6272 8730
rect 6324 8678 6336 8730
rect 6388 8678 6400 8730
rect 6452 8678 6464 8730
rect 6516 8678 9798 8730
rect 9850 8678 9862 8730
rect 9914 8678 9926 8730
rect 9978 8678 9990 8730
rect 10042 8678 11684 8730
rect 1104 8656 11684 8678
rect 3234 8616 3240 8628
rect 1872 8588 3240 8616
rect 1872 8412 1900 8588
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3418 8616 3424 8628
rect 3379 8588 3424 8616
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 9122 8616 9128 8628
rect 5040 8588 9128 8616
rect 5040 8576 5046 8588
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 9640 8588 10885 8616
rect 9640 8576 9646 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 4212 8520 6132 8548
rect 4212 8508 4218 8520
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 4430 8480 4436 8492
rect 2924 8452 3372 8480
rect 4391 8452 4436 8480
rect 2924 8440 2930 8452
rect 2133 8415 2191 8421
rect 2133 8412 2145 8415
rect 1872 8384 2145 8412
rect 2133 8381 2145 8384
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2332 8344 2360 8375
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 2639 8415 2697 8421
rect 2639 8412 2651 8415
rect 2464 8384 2651 8412
rect 2464 8372 2470 8384
rect 2639 8381 2651 8384
rect 2685 8381 2697 8415
rect 2639 8375 2697 8381
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 3050 8412 3056 8424
rect 2823 8384 3056 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3344 8421 3372 8452
rect 4430 8440 4436 8452
rect 4488 8480 4494 8492
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 4488 8452 5457 8480
rect 4488 8440 4494 8452
rect 5445 8449 5457 8452
rect 5491 8480 5503 8483
rect 6104 8480 6132 8520
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 7558 8548 7564 8560
rect 6880 8520 7564 8548
rect 6880 8508 6886 8520
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 5491 8452 5948 8480
rect 6104 8452 7941 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8381 3387 8415
rect 3602 8412 3608 8424
rect 3563 8384 3608 8412
rect 3329 8375 3387 8381
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 3881 8415 3939 8421
rect 3752 8384 3797 8412
rect 3752 8372 3758 8384
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 4338 8412 4344 8424
rect 4299 8384 4344 8412
rect 3881 8375 3939 8381
rect 2332 8316 2820 8344
rect 2792 8288 2820 8316
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3896 8344 3924 8375
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5074 8412 5080 8424
rect 5031 8384 5080 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 5258 8412 5264 8424
rect 5219 8384 5264 8412
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5920 8421 5948 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 7929 8443 7987 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8956 8452 9536 8480
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5408 8384 5549 8412
rect 5408 8372 5414 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 2924 8316 3924 8344
rect 5552 8344 5580 8375
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6052 8384 6377 8412
rect 6052 8372 6058 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 6687 8384 7297 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7466 8412 7472 8424
rect 7427 8384 7472 8412
rect 7285 8375 7343 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 7616 8384 7665 8412
rect 7616 8372 7622 8384
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 8956 8421 8984 8452
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8076 8384 8953 8412
rect 8076 8372 8082 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9122 8372 9128 8424
rect 9180 8412 9186 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 9180 8384 9229 8412
rect 9180 8372 9186 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9508 8412 9536 8452
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 9732 8452 10824 8480
rect 9732 8440 9738 8452
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 9508 8384 10057 8412
rect 9401 8375 9459 8381
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10318 8412 10324 8424
rect 10279 8384 10324 8412
rect 10045 8375 10103 8381
rect 6730 8344 6736 8356
rect 5552 8316 6736 8344
rect 2924 8304 2930 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 8294 8344 8300 8356
rect 6871 8316 8300 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 8389 8347 8447 8353
rect 8389 8313 8401 8347
rect 8435 8344 8447 8347
rect 9306 8344 9312 8356
rect 8435 8316 9312 8344
rect 8435 8313 8447 8316
rect 8389 8307 8447 8313
rect 1949 8279 2007 8285
rect 1949 8245 1961 8279
rect 1995 8276 2007 8279
rect 2682 8276 2688 8288
rect 1995 8248 2688 8276
rect 1995 8245 2007 8248
rect 1949 8239 2007 8245
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 5902 8276 5908 8288
rect 5500 8248 5908 8276
rect 5500 8236 5506 8248
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8404 8276 8432 8307
rect 9306 8304 9312 8316
rect 9364 8344 9370 8356
rect 9416 8344 9444 8375
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10686 8412 10692 8424
rect 10643 8384 10692 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 9364 8316 9444 8344
rect 9493 8347 9551 8353
rect 9364 8304 9370 8316
rect 9493 8313 9505 8347
rect 9539 8313 9551 8347
rect 10520 8344 10548 8375
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10796 8421 10824 8452
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 9493 8307 9551 8313
rect 10060 8316 10548 8344
rect 7892 8248 8432 8276
rect 7892 8236 7898 8248
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 9508 8276 9536 8307
rect 10060 8288 10088 8316
rect 10042 8276 10048 8288
rect 8904 8248 10048 8276
rect 8904 8236 8910 8248
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 1104 8186 11684 8208
rect 1104 8134 4508 8186
rect 4560 8134 4572 8186
rect 4624 8134 4636 8186
rect 4688 8134 4700 8186
rect 4752 8134 8035 8186
rect 8087 8134 8099 8186
rect 8151 8134 8163 8186
rect 8215 8134 8227 8186
rect 8279 8134 11684 8186
rect 1104 8112 11684 8134
rect 2148 8044 2636 8072
rect 2148 8013 2176 8044
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 7973 2191 8007
rect 2133 7967 2191 7973
rect 2498 7964 2504 8016
rect 2556 7964 2562 8016
rect 2608 8004 2636 8044
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2832 8044 2877 8072
rect 2832 8032 2838 8044
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 6178 8072 6184 8084
rect 3660 8044 6184 8072
rect 3660 8032 3666 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 7742 8072 7748 8084
rect 7576 8044 7748 8072
rect 3142 8004 3148 8016
rect 2608 7976 3148 8004
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 5353 8007 5411 8013
rect 5353 8004 5365 8007
rect 4356 7976 5365 8004
rect 2280 7939 2338 7945
rect 2280 7905 2292 7939
rect 2326 7936 2338 7939
rect 2516 7936 2544 7964
rect 4356 7945 4384 7976
rect 5353 7973 5365 7976
rect 5399 7973 5411 8007
rect 6914 8004 6920 8016
rect 5353 7967 5411 7973
rect 6104 7976 6920 8004
rect 2326 7908 2544 7936
rect 4341 7939 4399 7945
rect 2326 7905 2338 7908
rect 2280 7899 2338 7905
rect 4341 7905 4353 7939
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5810 7936 5816 7948
rect 5123 7908 5816 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 1452 7840 2513 7868
rect 1452 7828 1458 7840
rect 2501 7837 2513 7840
rect 2547 7868 2559 7871
rect 2682 7868 2688 7880
rect 2547 7840 2688 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 4430 7868 4436 7880
rect 4391 7840 4436 7868
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4816 7800 4844 7899
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6104 7945 6132 7976
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 7098 7936 7104 7948
rect 6319 7908 7104 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7466 7936 7472 7948
rect 7427 7908 7472 7936
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7576 7945 7604 8044
rect 7742 8032 7748 8044
rect 7800 8072 7806 8084
rect 8570 8072 8576 8084
rect 7800 8044 8576 8072
rect 7800 8032 7806 8044
rect 8570 8032 8576 8044
rect 8628 8072 8634 8084
rect 10962 8072 10968 8084
rect 8628 8044 9812 8072
rect 10923 8044 10968 8072
rect 8628 8032 8634 8044
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 7708 7976 7972 8004
rect 7708 7964 7714 7976
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 7944 7936 7972 7976
rect 8570 7936 8576 7948
rect 7883 7908 7972 7936
rect 8531 7908 8576 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 8720 7908 9689 7936
rect 8720 7896 8726 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9784 7936 9812 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 9907 7939 9965 7945
rect 9907 7936 9919 7939
rect 9784 7908 9919 7936
rect 9677 7899 9735 7905
rect 9907 7905 9919 7908
rect 9953 7905 9965 7939
rect 9907 7899 9965 7905
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10376 7908 10517 7936
rect 10376 7896 10382 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5994 7868 6000 7880
rect 5307 7840 6000 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7006 7868 7012 7880
rect 6963 7840 7012 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 6472 7800 6500 7831
rect 4816 7772 6500 7800
rect 6748 7800 6776 7831
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 8386 7868 8392 7880
rect 8343 7840 8392 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 8849 7871 8907 7877
rect 8849 7868 8861 7871
rect 8812 7840 8861 7868
rect 8812 7828 8818 7840
rect 8849 7837 8861 7840
rect 8895 7868 8907 7871
rect 9766 7868 9772 7880
rect 8895 7840 9772 7868
rect 8895 7837 8907 7840
rect 8849 7831 8907 7837
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10796 7868 10824 7899
rect 10336 7840 10824 7868
rect 10336 7812 10364 7840
rect 10137 7803 10195 7809
rect 10137 7800 10149 7803
rect 6748 7772 8432 7800
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7732 2470 7744
rect 3694 7732 3700 7744
rect 2464 7704 3700 7732
rect 2464 7692 2470 7704
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 6472 7732 6500 7772
rect 6730 7732 6736 7744
rect 6472 7704 6736 7732
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 8404 7732 8432 7772
rect 8588 7772 10149 7800
rect 8588 7732 8616 7772
rect 10137 7769 10149 7772
rect 10183 7769 10195 7803
rect 10137 7763 10195 7769
rect 10318 7760 10324 7812
rect 10376 7760 10382 7812
rect 8404 7704 8616 7732
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9815 7735 9873 7741
rect 9815 7732 9827 7735
rect 9364 7704 9827 7732
rect 9364 7692 9370 7704
rect 9815 7701 9827 7704
rect 9861 7701 9873 7735
rect 10594 7732 10600 7744
rect 10555 7704 10600 7732
rect 9815 7695 9873 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 1104 7642 11684 7664
rect 1104 7590 2745 7642
rect 2797 7590 2809 7642
rect 2861 7590 2873 7642
rect 2925 7590 2937 7642
rect 2989 7590 6272 7642
rect 6324 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 6464 7642
rect 6516 7590 9798 7642
rect 9850 7590 9862 7642
rect 9914 7590 9926 7642
rect 9978 7590 9990 7642
rect 10042 7590 11684 7642
rect 1104 7568 11684 7590
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7282 7528 7288 7540
rect 6963 7500 7288 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 8110 7528 8116 7540
rect 7524 7500 8116 7528
rect 7524 7488 7530 7500
rect 8110 7488 8116 7500
rect 8168 7528 8174 7540
rect 9582 7528 9588 7540
rect 8168 7500 9588 7528
rect 8168 7488 8174 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 5626 7460 5632 7472
rect 4264 7432 5632 7460
rect 4264 7333 4292 7432
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 6822 7460 6828 7472
rect 6380 7432 6828 7460
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 5353 7395 5411 7401
rect 4387 7364 4936 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4908 7336 4936 7364
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 6380 7392 6408 7432
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 8849 7463 8907 7469
rect 8849 7460 8861 7463
rect 7944 7432 8861 7460
rect 6638 7392 6644 7404
rect 5399 7364 6408 7392
rect 6472 7364 6644 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4706 7324 4712 7336
rect 4571 7296 4712 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4948 7296 4997 7324
rect 4948 7284 4954 7296
rect 4985 7293 4997 7296
rect 5031 7324 5043 7327
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5031 7296 5917 7324
rect 5031 7293 5043 7296
rect 4985 7287 5043 7293
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 6086 7324 6092 7336
rect 6047 7296 6092 7324
rect 5905 7287 5963 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 6472 7333 6500 7364
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6549 7287 6607 7293
rect 4617 7259 4675 7265
rect 4617 7225 4629 7259
rect 4663 7256 4675 7259
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4663 7228 4813 7256
rect 4663 7225 4675 7228
rect 4617 7219 4675 7225
rect 4801 7225 4813 7228
rect 4847 7256 4859 7259
rect 6564 7256 6592 7287
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 7944 7333 7972 7432
rect 8849 7429 8861 7432
rect 8895 7429 8907 7463
rect 8849 7423 8907 7429
rect 8938 7352 8944 7404
rect 8996 7392 9002 7404
rect 8996 7364 9904 7392
rect 8996 7352 9002 7364
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 8110 7324 8116 7336
rect 8071 7296 8116 7324
rect 7929 7287 7987 7293
rect 7190 7256 7196 7268
rect 4847 7228 6592 7256
rect 7151 7228 7196 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5000 7200 5028 7228
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 7760 7256 7788 7287
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8260 7296 8493 7324
rect 8260 7284 8266 7296
rect 8481 7293 8493 7296
rect 8527 7324 8539 7327
rect 8665 7327 8723 7333
rect 8527 7296 8616 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8386 7256 8392 7268
rect 7760 7228 8392 7256
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 4982 7148 4988 7200
rect 5040 7148 5046 7200
rect 5721 7191 5779 7197
rect 5721 7157 5733 7191
rect 5767 7188 5779 7191
rect 6914 7188 6920 7200
rect 5767 7160 6920 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 8588 7188 8616 7296
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8846 7324 8852 7336
rect 8807 7296 8852 7324
rect 8665 7287 8723 7293
rect 8680 7256 8708 7287
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 9582 7324 9588 7336
rect 9543 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9876 7333 9904 7364
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 10594 7256 10600 7268
rect 8680 7228 10600 7256
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 8588 7160 9689 7188
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9824 7160 9965 7188
rect 9824 7148 9830 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 1104 7098 11684 7120
rect 1104 7046 4508 7098
rect 4560 7046 4572 7098
rect 4624 7046 4636 7098
rect 4688 7046 4700 7098
rect 4752 7046 8035 7098
rect 8087 7046 8099 7098
rect 8151 7046 8163 7098
rect 8215 7046 8227 7098
rect 8279 7046 11684 7098
rect 1104 7024 11684 7046
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6822 6984 6828 6996
rect 5960 6956 6828 6984
rect 5960 6944 5966 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7558 6984 7564 6996
rect 7300 6956 7564 6984
rect 5442 6916 5448 6928
rect 5403 6888 5448 6916
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 7300 6916 7328 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9033 6987 9091 6993
rect 9033 6984 9045 6987
rect 8444 6956 9045 6984
rect 8444 6944 8450 6956
rect 9033 6953 9045 6956
rect 9079 6953 9091 6987
rect 9033 6947 9091 6953
rect 6052 6888 7328 6916
rect 6052 6876 6058 6888
rect 7742 6876 7748 6928
rect 7800 6916 7806 6928
rect 8846 6916 8852 6928
rect 7800 6888 8156 6916
rect 7800 6876 7806 6888
rect 4890 6848 4896 6860
rect 4851 6820 4896 6848
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5040 6820 5085 6848
rect 5040 6808 5046 6820
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 6086 6848 6092 6860
rect 5960 6820 6092 6848
rect 5960 6808 5966 6820
rect 6086 6808 6092 6820
rect 6144 6848 6150 6860
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 6144 6820 6193 6848
rect 6144 6808 6150 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6638 6848 6644 6860
rect 6595 6820 6644 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7616 6820 7665 6848
rect 7616 6808 7622 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7926 6848 7932 6860
rect 7653 6811 7711 6817
rect 7760 6820 7932 6848
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5684 6752 6009 6780
rect 5684 6740 5690 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 7377 6783 7435 6789
rect 6871 6752 7328 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 5534 6712 5540 6724
rect 4856 6684 5540 6712
rect 4856 6672 4862 6684
rect 5534 6672 5540 6684
rect 5592 6712 5598 6724
rect 6178 6712 6184 6724
rect 5592 6684 6184 6712
rect 5592 6672 5598 6684
rect 6178 6672 6184 6684
rect 6236 6712 6242 6724
rect 6472 6712 6500 6743
rect 6236 6684 6500 6712
rect 6236 6672 6242 6684
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 6086 6644 6092 6656
rect 5859 6616 6092 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 7300 6644 7328 6752
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7760 6780 7788 6820
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 7423 6752 7788 6780
rect 7837 6783 7895 6789
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 8128 6780 8156 6888
rect 8312 6888 8852 6916
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8312 6848 8340 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 10318 6916 10324 6928
rect 9732 6888 10324 6916
rect 9732 6876 9738 6888
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 8251 6820 8340 6848
rect 8389 6851 8447 6857
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8389 6817 8401 6851
rect 8435 6817 8447 6851
rect 8757 6851 8815 6857
rect 8757 6848 8769 6851
rect 8389 6811 8447 6817
rect 8588 6820 8769 6848
rect 8404 6780 8432 6811
rect 8588 6792 8616 6820
rect 8757 6817 8769 6820
rect 8803 6817 8815 6851
rect 8938 6848 8944 6860
rect 8899 6820 8944 6848
rect 8757 6811 8815 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10686 6848 10692 6860
rect 9907 6820 10692 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 8570 6780 8576 6792
rect 8128 6752 8432 6780
rect 8531 6752 8576 6780
rect 7837 6743 7895 6749
rect 7650 6644 7656 6656
rect 7300 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6644 7714 6656
rect 7852 6644 7880 6743
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8662 6644 8668 6656
rect 7708 6616 8668 6644
rect 7708 6604 7714 6616
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10134 6644 10140 6656
rect 9999 6616 10140 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 1104 6554 11684 6576
rect 1104 6502 2745 6554
rect 2797 6502 2809 6554
rect 2861 6502 2873 6554
rect 2925 6502 2937 6554
rect 2989 6502 6272 6554
rect 6324 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 6464 6554
rect 6516 6502 9798 6554
rect 9850 6502 9862 6554
rect 9914 6502 9926 6554
rect 9978 6502 9990 6554
rect 10042 6502 11684 6554
rect 1104 6480 11684 6502
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 6638 6440 6644 6452
rect 5951 6412 6644 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7156 6412 7941 6440
rect 7156 6400 7162 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 10686 6440 10692 6452
rect 10647 6412 10692 6440
rect 7929 6403 7987 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 9674 6372 9680 6384
rect 6840 6344 9680 6372
rect 5810 6264 5816 6316
rect 5868 6304 5874 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 5868 6276 6561 6304
rect 5868 6264 5874 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 3292 6208 5641 6236
rect 3292 6196 3298 6208
rect 5629 6205 5641 6208
rect 5675 6236 5687 6239
rect 5718 6236 5724 6248
rect 5675 6208 5724 6236
rect 5675 6205 5687 6208
rect 5629 6199 5687 6205
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 6086 6236 6092 6248
rect 6047 6208 6092 6236
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 6270 6236 6276 6248
rect 6183 6208 6276 6236
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 6840 6245 6868 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10410 6372 10416 6384
rect 9824 6344 10416 6372
rect 9824 6332 9830 6344
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 7484 6276 8401 6304
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7374 6236 7380 6248
rect 7147 6208 7380 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 2406 6128 2412 6180
rect 2464 6168 2470 6180
rect 6288 6168 6316 6196
rect 2464 6140 6316 6168
rect 6932 6168 6960 6199
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7282 6168 7288 6180
rect 6932 6140 7288 6168
rect 2464 6128 2470 6140
rect 7282 6128 7288 6140
rect 7340 6128 7346 6180
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7484 6100 7512 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 9306 6304 9312 6316
rect 8389 6267 8447 6273
rect 8496 6276 9312 6304
rect 7650 6236 7656 6248
rect 7611 6208 7656 6236
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 7834 6236 7840 6248
rect 7795 6208 7840 6236
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6236 8355 6239
rect 8496 6236 8524 6276
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 8343 6208 8524 6236
rect 9125 6239 9183 6245
rect 8343 6205 8355 6208
rect 8297 6199 8355 6205
rect 9125 6205 9137 6239
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 7561 6171 7619 6177
rect 7561 6137 7573 6171
rect 7607 6137 7619 6171
rect 7561 6131 7619 6137
rect 6788 6072 7512 6100
rect 7576 6100 7604 6131
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 9140 6168 9168 6199
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9677 6239 9735 6245
rect 9272 6208 9317 6236
rect 9272 6196 9278 6208
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 9766 6236 9772 6248
rect 9723 6208 9772 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6236 9919 6239
rect 10134 6236 10140 6248
rect 9907 6208 10140 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 9876 6168 9904 6199
rect 10134 6196 10140 6208
rect 10192 6236 10198 6248
rect 10192 6208 10272 6236
rect 10192 6196 10198 6208
rect 7800 6140 9076 6168
rect 9140 6140 9904 6168
rect 7800 6128 7806 6140
rect 7834 6100 7840 6112
rect 7576 6072 7840 6100
rect 6788 6060 6794 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 9048 6100 9076 6140
rect 9122 6100 9128 6112
rect 9048 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9732 6072 10149 6100
rect 9732 6060 9738 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10244 6100 10272 6208
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 10376 6208 10425 6236
rect 10376 6196 10382 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10594 6236 10600 6248
rect 10555 6208 10600 6236
rect 10413 6199 10471 6205
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 10594 6100 10600 6112
rect 10244 6072 10600 6100
rect 10137 6063 10195 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 1104 6010 11684 6032
rect 1104 5958 4508 6010
rect 4560 5958 4572 6010
rect 4624 5958 4636 6010
rect 4688 5958 4700 6010
rect 4752 5958 8035 6010
rect 8087 5958 8099 6010
rect 8151 5958 8163 6010
rect 8215 5958 8227 6010
rect 8279 5958 11684 6010
rect 1104 5936 11684 5958
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 5960 5868 6377 5896
rect 5960 5856 5966 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 8938 5896 8944 5908
rect 7699 5868 8944 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 10686 5856 10692 5908
rect 10744 5856 10750 5908
rect 7469 5831 7527 5837
rect 7469 5797 7481 5831
rect 7515 5828 7527 5831
rect 7742 5828 7748 5840
rect 7515 5800 7748 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 7926 5828 7932 5840
rect 7887 5800 7932 5828
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 10704 5828 10732 5856
rect 10336 5800 10732 5828
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 3200 5732 6285 5760
rect 3200 5720 3206 5732
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 6273 5723 6331 5729
rect 6288 5692 6316 5723
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7193 5763 7251 5769
rect 7193 5760 7205 5763
rect 6972 5732 7205 5760
rect 6972 5720 6978 5732
rect 7193 5729 7205 5732
rect 7239 5729 7251 5763
rect 7193 5723 7251 5729
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 7650 5760 7656 5772
rect 7607 5732 7656 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7834 5760 7840 5772
rect 7795 5732 7840 5760
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 10336 5769 10364 5800
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5760 10747 5763
rect 10778 5760 10784 5772
rect 10735 5732 10784 5760
rect 10735 5729 10747 5732
rect 10689 5723 10747 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 6288 5664 9689 5692
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 9677 5655 9735 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10594 5692 10600 5704
rect 10555 5664 10600 5692
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 7282 5584 7288 5636
rect 7340 5624 7346 5636
rect 8570 5624 8576 5636
rect 7340 5596 8576 5624
rect 7340 5584 7346 5596
rect 8570 5584 8576 5596
rect 8628 5624 8634 5636
rect 9030 5624 9036 5636
rect 8628 5596 9036 5624
rect 8628 5584 8634 5596
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 9674 5556 9680 5568
rect 5776 5528 9680 5556
rect 5776 5516 5782 5528
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 1104 5466 11684 5488
rect 1104 5414 2745 5466
rect 2797 5414 2809 5466
rect 2861 5414 2873 5466
rect 2925 5414 2937 5466
rect 2989 5414 6272 5466
rect 6324 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 6464 5466
rect 6516 5414 9798 5466
rect 9850 5414 9862 5466
rect 9914 5414 9926 5466
rect 9978 5414 9990 5466
rect 10042 5414 11684 5466
rect 1104 5392 11684 5414
rect 1104 4922 11684 4944
rect 1104 4870 4508 4922
rect 4560 4870 4572 4922
rect 4624 4870 4636 4922
rect 4688 4870 4700 4922
rect 4752 4870 8035 4922
rect 8087 4870 8099 4922
rect 8151 4870 8163 4922
rect 8215 4870 8227 4922
rect 8279 4870 11684 4922
rect 1104 4848 11684 4870
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 474 4428 480 4480
rect 532 4468 538 4480
rect 1581 4471 1639 4477
rect 1581 4468 1593 4471
rect 532 4440 1593 4468
rect 532 4428 538 4440
rect 1581 4437 1593 4440
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 1104 4378 11684 4400
rect 1104 4326 2745 4378
rect 2797 4326 2809 4378
rect 2861 4326 2873 4378
rect 2925 4326 2937 4378
rect 2989 4326 6272 4378
rect 6324 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 6464 4378
rect 6516 4326 9798 4378
rect 9850 4326 9862 4378
rect 9914 4326 9926 4378
rect 9978 4326 9990 4378
rect 10042 4326 11684 4378
rect 1104 4304 11684 4326
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5626 4128 5632 4140
rect 4856 4100 5632 4128
rect 4856 4088 4862 4100
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 1104 3834 11684 3856
rect 1104 3782 4508 3834
rect 4560 3782 4572 3834
rect 4624 3782 4636 3834
rect 4688 3782 4700 3834
rect 4752 3782 8035 3834
rect 8087 3782 8099 3834
rect 8151 3782 8163 3834
rect 8215 3782 8227 3834
rect 8279 3782 11684 3834
rect 1104 3760 11684 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 6822 3720 6828 3732
rect 2648 3692 6828 3720
rect 2648 3680 2654 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10560 3692 10885 3720
rect 10560 3680 10566 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 7248 3624 10456 3652
rect 7248 3612 7254 3624
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3584 9919 3587
rect 10226 3584 10232 3596
rect 9907 3556 10232 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 10226 3544 10232 3556
rect 10284 3584 10290 3596
rect 10428 3593 10456 3624
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 10284 3556 10333 3584
rect 10284 3544 10290 3556
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 9784 3448 9812 3479
rect 12158 3448 12164 3460
rect 9784 3420 12164 3448
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 1104 3290 11684 3312
rect 1104 3238 2745 3290
rect 2797 3238 2809 3290
rect 2861 3238 2873 3290
rect 2925 3238 2937 3290
rect 2989 3238 6272 3290
rect 6324 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 6464 3290
rect 6516 3238 9798 3290
rect 9850 3238 9862 3290
rect 9914 3238 9926 3290
rect 9978 3238 9990 3290
rect 10042 3238 11684 3290
rect 1104 3216 11684 3238
rect 10226 3176 10232 3188
rect 10187 3148 10232 3176
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 9125 3111 9183 3117
rect 9125 3077 9137 3111
rect 9171 3108 9183 3111
rect 10134 3108 10140 3120
rect 9171 3080 10140 3108
rect 9171 3077 9183 3080
rect 9125 3071 9183 3077
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 10244 3040 10272 3136
rect 7064 3012 9904 3040
rect 7064 3000 7070 3012
rect 9876 2981 9904 3012
rect 9968 3012 10272 3040
rect 9968 2981 9996 3012
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 9309 2935 9367 2941
rect 9493 2975 9551 2981
rect 9493 2941 9505 2975
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 9953 2975 10011 2981
rect 9953 2941 9965 2975
rect 9999 2941 10011 2975
rect 10134 2972 10140 2984
rect 10095 2944 10140 2972
rect 9953 2935 10011 2941
rect 9324 2836 9352 2935
rect 9508 2904 9536 2935
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 10152 2904 10180 2932
rect 9508 2876 10180 2904
rect 11054 2836 11060 2848
rect 9324 2808 11060 2836
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 1104 2746 11684 2768
rect 1104 2694 4508 2746
rect 4560 2694 4572 2746
rect 4624 2694 4636 2746
rect 4688 2694 4700 2746
rect 4752 2694 8035 2746
rect 8087 2694 8099 2746
rect 8151 2694 8163 2746
rect 8215 2694 8227 2746
rect 8279 2694 11684 2746
rect 1104 2672 11684 2694
rect 10045 2635 10103 2641
rect 10045 2601 10057 2635
rect 10091 2632 10103 2635
rect 10134 2632 10140 2644
rect 10091 2604 10140 2632
rect 10091 2601 10103 2604
rect 10045 2595 10103 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 8205 2499 8263 2505
rect 8205 2496 8217 2499
rect 7248 2468 8217 2496
rect 7248 2456 7254 2468
rect 8205 2465 8217 2468
rect 8251 2465 8263 2499
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 8205 2459 8263 2465
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 8628 2468 9781 2496
rect 8628 2456 8634 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 10134 2496 10140 2508
rect 9999 2468 10140 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 7984 2264 8309 2292
rect 7984 2252 7990 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 8757 2295 8815 2301
rect 8757 2261 8769 2295
rect 8803 2292 8815 2295
rect 8938 2292 8944 2304
rect 8803 2264 8944 2292
rect 8803 2261 8815 2264
rect 8757 2255 8815 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 1104 2202 11684 2224
rect 1104 2150 2745 2202
rect 2797 2150 2809 2202
rect 2861 2150 2873 2202
rect 2925 2150 2937 2202
rect 2989 2150 6272 2202
rect 6324 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 6464 2202
rect 6516 2150 9798 2202
rect 9850 2150 9862 2202
rect 9914 2150 9926 2202
rect 9978 2150 9990 2202
rect 10042 2150 11684 2202
rect 1104 2128 11684 2150
<< via1 >>
rect 4508 12486 4560 12538
rect 4572 12486 4624 12538
rect 4636 12486 4688 12538
rect 4700 12486 4752 12538
rect 8035 12486 8087 12538
rect 8099 12486 8151 12538
rect 8163 12486 8215 12538
rect 8227 12486 8279 12538
rect 5724 12248 5776 12300
rect 8944 12248 8996 12300
rect 4068 12180 4120 12232
rect 5448 12044 5500 12096
rect 7656 12044 7708 12096
rect 2745 11942 2797 11994
rect 2809 11942 2861 11994
rect 2873 11942 2925 11994
rect 2937 11942 2989 11994
rect 6272 11942 6324 11994
rect 6336 11942 6388 11994
rect 6400 11942 6452 11994
rect 6464 11942 6516 11994
rect 9798 11942 9850 11994
rect 9862 11942 9914 11994
rect 9926 11942 9978 11994
rect 9990 11942 10042 11994
rect 1492 11704 1544 11756
rect 1860 11704 1912 11756
rect 2780 11636 2832 11688
rect 3608 11704 3660 11756
rect 7932 11704 7984 11756
rect 4068 11636 4120 11688
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 7932 11568 7984 11620
rect 5724 11500 5776 11552
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 4508 11398 4560 11450
rect 4572 11398 4624 11450
rect 4636 11398 4688 11450
rect 4700 11398 4752 11450
rect 8035 11398 8087 11450
rect 8099 11398 8151 11450
rect 8163 11398 8215 11450
rect 8227 11398 8279 11450
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 7012 11228 7064 11280
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4804 11160 4856 11212
rect 6092 11160 6144 11212
rect 7656 11203 7708 11212
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 10416 11160 10468 11212
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 5540 11092 5592 11101
rect 480 11024 532 11076
rect 1492 11024 1544 11076
rect 8392 11092 8444 11144
rect 8300 11024 8352 11076
rect 6828 10956 6880 11008
rect 2745 10854 2797 10906
rect 2809 10854 2861 10906
rect 2873 10854 2925 10906
rect 2937 10854 2989 10906
rect 6272 10854 6324 10906
rect 6336 10854 6388 10906
rect 6400 10854 6452 10906
rect 6464 10854 6516 10906
rect 9798 10854 9850 10906
rect 9862 10854 9914 10906
rect 9926 10854 9978 10906
rect 9990 10854 10042 10906
rect 7656 10752 7708 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 6000 10684 6052 10736
rect 5632 10616 5684 10668
rect 5816 10548 5868 10600
rect 8852 10684 8904 10736
rect 9680 10684 9732 10736
rect 7748 10616 7800 10668
rect 7840 10616 7892 10668
rect 4896 10480 4948 10532
rect 6644 10548 6696 10600
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 8760 10548 8812 10600
rect 6920 10480 6972 10532
rect 8392 10480 8444 10532
rect 9036 10480 9088 10532
rect 6828 10412 6880 10464
rect 9680 10412 9732 10464
rect 4508 10310 4560 10362
rect 4572 10310 4624 10362
rect 4636 10310 4688 10362
rect 4700 10310 4752 10362
rect 8035 10310 8087 10362
rect 8099 10310 8151 10362
rect 8163 10310 8215 10362
rect 8227 10310 8279 10362
rect 5080 10208 5132 10260
rect 5816 10208 5868 10260
rect 4068 10140 4120 10192
rect 5632 10140 5684 10192
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 4344 10072 4396 10124
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 3056 10004 3108 10056
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 5816 10072 5868 10124
rect 6736 10072 6788 10124
rect 8668 10208 8720 10260
rect 7472 10140 7524 10192
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 8392 10072 8444 10124
rect 8852 10072 8904 10124
rect 7012 10004 7064 10056
rect 3424 9936 3476 9988
rect 4804 9936 4856 9988
rect 5632 9936 5684 9988
rect 9404 10004 9456 10056
rect 8484 9936 8536 9988
rect 7656 9868 7708 9920
rect 7932 9868 7984 9920
rect 8944 9868 8996 9920
rect 9128 9868 9180 9920
rect 2745 9766 2797 9818
rect 2809 9766 2861 9818
rect 2873 9766 2925 9818
rect 2937 9766 2989 9818
rect 6272 9766 6324 9818
rect 6336 9766 6388 9818
rect 6400 9766 6452 9818
rect 6464 9766 6516 9818
rect 9798 9766 9850 9818
rect 9862 9766 9914 9818
rect 9926 9766 9978 9818
rect 9990 9766 10042 9818
rect 3700 9664 3752 9716
rect 5264 9664 5316 9716
rect 5448 9664 5500 9716
rect 7288 9664 7340 9716
rect 7932 9664 7984 9716
rect 10324 9664 10376 9716
rect 10508 9664 10560 9716
rect 12164 9664 12216 9716
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 4988 9460 5040 9512
rect 5448 9460 5500 9512
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 6092 9528 6144 9580
rect 2412 9324 2464 9376
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8576 9528 8628 9580
rect 6920 9460 6972 9512
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7932 9460 7984 9512
rect 9036 9460 9088 9512
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 10692 9596 10744 9648
rect 9496 9528 9548 9580
rect 10232 9460 10284 9512
rect 11060 9460 11112 9512
rect 5356 9324 5408 9376
rect 5724 9324 5776 9376
rect 6276 9324 6328 9376
rect 9496 9392 9548 9444
rect 10600 9324 10652 9376
rect 4508 9222 4560 9274
rect 4572 9222 4624 9274
rect 4636 9222 4688 9274
rect 4700 9222 4752 9274
rect 8035 9222 8087 9274
rect 8099 9222 8151 9274
rect 8163 9222 8215 9274
rect 8227 9222 8279 9274
rect 2504 9120 2556 9172
rect 5816 9120 5868 9172
rect 6184 9120 6236 9172
rect 6828 9120 6880 9172
rect 7288 9120 7340 9172
rect 9220 9120 9272 9172
rect 9496 9120 9548 9172
rect 10600 9163 10652 9172
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 3056 8984 3108 9036
rect 3700 9027 3752 9036
rect 3700 8993 3709 9027
rect 3709 8993 3743 9027
rect 3743 8993 3752 9027
rect 3700 8984 3752 8993
rect 5172 9052 5224 9104
rect 5264 9052 5316 9104
rect 10600 9129 10609 9163
rect 10609 9129 10643 9163
rect 10643 9129 10652 9163
rect 10600 9120 10652 9129
rect 10784 9120 10836 9172
rect 4436 8984 4488 9036
rect 5448 8984 5500 9036
rect 6276 8984 6328 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7012 9027 7064 9036
rect 7012 8993 7021 9027
rect 7021 8993 7055 9027
rect 7055 8993 7064 9027
rect 7012 8984 7064 8993
rect 8760 9027 8812 9036
rect 5816 8916 5868 8968
rect 6184 8916 6236 8968
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 6736 8916 6788 8968
rect 7012 8848 7064 8900
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 8760 8984 8812 8993
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9772 8984 9824 9036
rect 10508 9027 10560 9036
rect 8208 8848 8260 8900
rect 9128 8916 9180 8968
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 8668 8848 8720 8900
rect 1492 8780 1544 8832
rect 3608 8780 3660 8832
rect 7472 8780 7524 8832
rect 7564 8780 7616 8832
rect 8852 8780 8904 8832
rect 9036 8780 9088 8832
rect 9312 8780 9364 8832
rect 2745 8678 2797 8730
rect 2809 8678 2861 8730
rect 2873 8678 2925 8730
rect 2937 8678 2989 8730
rect 6272 8678 6324 8730
rect 6336 8678 6388 8730
rect 6400 8678 6452 8730
rect 6464 8678 6516 8730
rect 9798 8678 9850 8730
rect 9862 8678 9914 8730
rect 9926 8678 9978 8730
rect 9990 8678 10042 8730
rect 3240 8576 3292 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 4988 8576 5040 8628
rect 9128 8576 9180 8628
rect 9588 8576 9640 8628
rect 4160 8508 4212 8560
rect 2872 8440 2924 8492
rect 4436 8483 4488 8492
rect 2412 8372 2464 8424
rect 3056 8372 3108 8424
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 6828 8508 6880 8560
rect 7564 8508 7616 8560
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 4344 8415 4396 8424
rect 2872 8304 2924 8356
rect 4344 8381 4353 8415
rect 4353 8381 4387 8415
rect 4387 8381 4396 8415
rect 4344 8372 4396 8381
rect 5080 8372 5132 8424
rect 5264 8415 5316 8424
rect 5264 8381 5273 8415
rect 5273 8381 5307 8415
rect 5307 8381 5316 8415
rect 5264 8372 5316 8381
rect 5356 8372 5408 8424
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 6000 8372 6052 8424
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 7564 8372 7616 8424
rect 8024 8372 8076 8424
rect 9128 8372 9180 8424
rect 9680 8440 9732 8492
rect 10324 8415 10376 8424
rect 6736 8304 6788 8356
rect 8300 8304 8352 8356
rect 2688 8236 2740 8288
rect 2780 8236 2832 8288
rect 5448 8236 5500 8288
rect 5908 8236 5960 8288
rect 7840 8236 7892 8288
rect 9312 8304 9364 8356
rect 10324 8381 10333 8415
rect 10333 8381 10367 8415
rect 10367 8381 10376 8415
rect 10324 8372 10376 8381
rect 10692 8372 10744 8424
rect 8852 8236 8904 8288
rect 10048 8236 10100 8288
rect 4508 8134 4560 8186
rect 4572 8134 4624 8186
rect 4636 8134 4688 8186
rect 4700 8134 4752 8186
rect 8035 8134 8087 8186
rect 8099 8134 8151 8186
rect 8163 8134 8215 8186
rect 8227 8134 8279 8186
rect 2504 7964 2556 8016
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 3608 8032 3660 8084
rect 6184 8032 6236 8084
rect 3148 7964 3200 8016
rect 5816 7939 5868 7948
rect 1400 7828 1452 7880
rect 2688 7828 2740 7880
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6920 7964 6972 8016
rect 7104 7896 7156 7948
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 7748 8032 7800 8084
rect 8576 8032 8628 8084
rect 10968 8075 11020 8084
rect 7656 7964 7708 8016
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 8668 7896 8720 7948
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 10324 7896 10376 7948
rect 6000 7828 6052 7880
rect 7012 7828 7064 7880
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8392 7828 8444 7880
rect 8760 7828 8812 7880
rect 9772 7828 9824 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3700 7692 3752 7744
rect 6736 7692 6788 7744
rect 10324 7760 10376 7812
rect 9312 7692 9364 7744
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 2745 7590 2797 7642
rect 2809 7590 2861 7642
rect 2873 7590 2925 7642
rect 2937 7590 2989 7642
rect 6272 7590 6324 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 6464 7590 6516 7642
rect 9798 7590 9850 7642
rect 9862 7590 9914 7642
rect 9926 7590 9978 7642
rect 9990 7590 10042 7642
rect 7288 7488 7340 7540
rect 7472 7488 7524 7540
rect 8116 7488 8168 7540
rect 9588 7488 9640 7540
rect 5632 7420 5684 7472
rect 6828 7420 6880 7472
rect 4712 7284 4764 7336
rect 4896 7284 4948 7336
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 6644 7352 6696 7404
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8944 7352 8996 7404
rect 8116 7327 8168 7336
rect 7196 7259 7248 7268
rect 7196 7225 7205 7259
rect 7205 7225 7239 7259
rect 7239 7225 7248 7259
rect 7196 7216 7248 7225
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 8208 7284 8260 7336
rect 8392 7216 8444 7268
rect 4988 7148 5040 7200
rect 6920 7148 6972 7200
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 10600 7216 10652 7268
rect 9772 7148 9824 7200
rect 4508 7046 4560 7098
rect 4572 7046 4624 7098
rect 4636 7046 4688 7098
rect 4700 7046 4752 7098
rect 8035 7046 8087 7098
rect 8099 7046 8151 7098
rect 8163 7046 8215 7098
rect 8227 7046 8279 7098
rect 5908 6944 5960 6996
rect 6828 6944 6880 6996
rect 5448 6919 5500 6928
rect 5448 6885 5457 6919
rect 5457 6885 5491 6919
rect 5491 6885 5500 6919
rect 5448 6876 5500 6885
rect 6000 6876 6052 6928
rect 7564 6944 7616 6996
rect 8392 6944 8444 6996
rect 7748 6876 7800 6928
rect 4896 6851 4948 6860
rect 4896 6817 4905 6851
rect 4905 6817 4939 6851
rect 4939 6817 4948 6851
rect 4896 6808 4948 6817
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5908 6808 5960 6860
rect 6092 6808 6144 6860
rect 6644 6808 6696 6860
rect 7564 6808 7616 6860
rect 5632 6740 5684 6792
rect 4804 6672 4856 6724
rect 5540 6672 5592 6724
rect 6184 6672 6236 6724
rect 6092 6604 6144 6656
rect 7932 6808 7984 6860
rect 8852 6876 8904 6928
rect 9680 6876 9732 6928
rect 10324 6876 10376 6928
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 10692 6808 10744 6860
rect 8576 6783 8628 6792
rect 7656 6604 7708 6656
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8668 6604 8720 6656
rect 10140 6604 10192 6656
rect 2745 6502 2797 6554
rect 2809 6502 2861 6554
rect 2873 6502 2925 6554
rect 2937 6502 2989 6554
rect 6272 6502 6324 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 6464 6502 6516 6554
rect 9798 6502 9850 6554
rect 9862 6502 9914 6554
rect 9926 6502 9978 6554
rect 9990 6502 10042 6554
rect 6644 6400 6696 6452
rect 7104 6400 7156 6452
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 5816 6264 5868 6316
rect 3240 6196 3292 6248
rect 5724 6196 5776 6248
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 6276 6239 6328 6248
rect 6276 6205 6285 6239
rect 6285 6205 6319 6239
rect 6319 6205 6328 6239
rect 6276 6196 6328 6205
rect 9680 6332 9732 6384
rect 9772 6332 9824 6384
rect 10416 6332 10468 6384
rect 2412 6128 2464 6180
rect 7380 6196 7432 6248
rect 7288 6128 7340 6180
rect 6736 6060 6788 6112
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 9312 6264 9364 6316
rect 7748 6128 7800 6180
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 9772 6196 9824 6248
rect 10140 6196 10192 6248
rect 7840 6060 7892 6112
rect 9128 6060 9180 6112
rect 9680 6060 9732 6112
rect 10324 6196 10376 6248
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 10600 6060 10652 6112
rect 4508 5958 4560 6010
rect 4572 5958 4624 6010
rect 4636 5958 4688 6010
rect 4700 5958 4752 6010
rect 8035 5958 8087 6010
rect 8099 5958 8151 6010
rect 8163 5958 8215 6010
rect 8227 5958 8279 6010
rect 5908 5856 5960 5908
rect 8944 5856 8996 5908
rect 10692 5856 10744 5908
rect 7748 5788 7800 5840
rect 7932 5831 7984 5840
rect 7932 5797 7941 5831
rect 7941 5797 7975 5831
rect 7975 5797 7984 5831
rect 7932 5788 7984 5797
rect 3148 5720 3200 5772
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 6920 5720 6972 5772
rect 7656 5720 7708 5772
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 10784 5720 10836 5772
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 7288 5584 7340 5636
rect 8576 5584 8628 5636
rect 9036 5584 9088 5636
rect 5724 5516 5776 5568
rect 9680 5516 9732 5568
rect 2745 5414 2797 5466
rect 2809 5414 2861 5466
rect 2873 5414 2925 5466
rect 2937 5414 2989 5466
rect 6272 5414 6324 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 6464 5414 6516 5466
rect 9798 5414 9850 5466
rect 9862 5414 9914 5466
rect 9926 5414 9978 5466
rect 9990 5414 10042 5466
rect 4508 4870 4560 4922
rect 4572 4870 4624 4922
rect 4636 4870 4688 4922
rect 4700 4870 4752 4922
rect 8035 4870 8087 4922
rect 8099 4870 8151 4922
rect 8163 4870 8215 4922
rect 8227 4870 8279 4922
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 480 4428 532 4480
rect 2745 4326 2797 4378
rect 2809 4326 2861 4378
rect 2873 4326 2925 4378
rect 2937 4326 2989 4378
rect 6272 4326 6324 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 6464 4326 6516 4378
rect 9798 4326 9850 4378
rect 9862 4326 9914 4378
rect 9926 4326 9978 4378
rect 9990 4326 10042 4378
rect 4804 4088 4856 4140
rect 5632 4088 5684 4140
rect 4508 3782 4560 3834
rect 4572 3782 4624 3834
rect 4636 3782 4688 3834
rect 4700 3782 4752 3834
rect 8035 3782 8087 3834
rect 8099 3782 8151 3834
rect 8163 3782 8215 3834
rect 8227 3782 8279 3834
rect 2596 3680 2648 3732
rect 6828 3680 6880 3732
rect 10508 3680 10560 3732
rect 7196 3612 7248 3664
rect 10232 3544 10284 3596
rect 12164 3408 12216 3460
rect 2745 3238 2797 3290
rect 2809 3238 2861 3290
rect 2873 3238 2925 3290
rect 2937 3238 2989 3290
rect 6272 3238 6324 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 6464 3238 6516 3290
rect 9798 3238 9850 3290
rect 9862 3238 9914 3290
rect 9926 3238 9978 3290
rect 9990 3238 10042 3290
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 10140 3068 10192 3120
rect 7012 3000 7064 3052
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 11060 2796 11112 2848
rect 4508 2694 4560 2746
rect 4572 2694 4624 2746
rect 4636 2694 4688 2746
rect 4700 2694 4752 2746
rect 8035 2694 8087 2746
rect 8099 2694 8151 2746
rect 8163 2694 8215 2746
rect 8227 2694 8279 2746
rect 10140 2592 10192 2644
rect 7196 2456 7248 2508
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 10140 2456 10192 2508
rect 7932 2252 7984 2304
rect 8944 2252 8996 2304
rect 2745 2150 2797 2202
rect 2809 2150 2861 2202
rect 2873 2150 2925 2202
rect 2937 2150 2989 2202
rect 6272 2150 6324 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
rect 6464 2150 6516 2202
rect 9798 2150 9850 2202
rect 9862 2150 9914 2202
rect 9926 2150 9978 2202
rect 9990 2150 10042 2202
<< metal2 >>
rect 478 14167 534 14967
rect 1490 14167 1546 14967
rect 2594 14167 2650 14967
rect 3606 14167 3662 14967
rect 4710 14167 4766 14967
rect 5722 14167 5778 14967
rect 6826 14167 6882 14967
rect 7930 14167 7986 14967
rect 8942 14167 8998 14967
rect 10046 14167 10102 14967
rect 11058 14167 11114 14967
rect 12162 14167 12218 14967
rect 492 11082 520 14167
rect 1504 11762 1532 14167
rect 2608 11778 2636 14167
rect 3054 13696 3110 13705
rect 3054 13631 3110 13640
rect 2719 11996 3015 12016
rect 2775 11994 2799 11996
rect 2855 11994 2879 11996
rect 2935 11994 2959 11996
rect 2797 11942 2799 11994
rect 2861 11942 2873 11994
rect 2935 11942 2937 11994
rect 2775 11940 2799 11942
rect 2855 11940 2879 11942
rect 2935 11940 2959 11942
rect 2719 11920 3015 11940
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1860 11756 1912 11762
rect 2608 11750 2820 11778
rect 1860 11698 1912 11704
rect 1398 11248 1454 11257
rect 1398 11183 1454 11192
rect 480 11076 532 11082
rect 480 11018 532 11024
rect 1412 9518 1440 11183
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1504 10033 1532 11018
rect 1490 10024 1546 10033
rect 1490 9959 1546 9968
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1504 9330 1532 9959
rect 1412 9302 1532 9330
rect 1412 7886 1440 9302
rect 1872 9042 1900 11698
rect 2792 11694 2820 11750
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2719 10908 3015 10928
rect 2775 10906 2799 10908
rect 2855 10906 2879 10908
rect 2935 10906 2959 10908
rect 2797 10854 2799 10906
rect 2861 10854 2873 10906
rect 2935 10854 2937 10906
rect 2775 10852 2799 10854
rect 2855 10852 2879 10854
rect 2935 10852 2959 10854
rect 2719 10832 3015 10852
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 1492 8832 1544 8838
rect 2240 8809 2268 8978
rect 1492 8774 1544 8780
rect 2226 8800 2282 8809
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 4690 1440 7822
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 480 4480 532 4486
rect 480 4422 532 4428
rect 492 800 520 4422
rect 1504 800 1532 8774
rect 2226 8735 2282 8744
rect 2424 8430 2452 9318
rect 2516 9178 2544 10066
rect 3068 10062 3096 13631
rect 3620 11762 3648 14167
rect 4724 12730 4752 14167
rect 4724 12702 4844 12730
rect 4482 12540 4778 12560
rect 4538 12538 4562 12540
rect 4618 12538 4642 12540
rect 4698 12538 4722 12540
rect 4560 12486 4562 12538
rect 4624 12486 4636 12538
rect 4698 12486 4700 12538
rect 4538 12484 4562 12486
rect 4618 12484 4642 12486
rect 4698 12484 4722 12486
rect 4482 12464 4778 12484
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 4080 11694 4108 12174
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11218 4108 11630
rect 4482 11452 4778 11472
rect 4538 11450 4562 11452
rect 4618 11450 4642 11452
rect 4698 11450 4722 11452
rect 4560 11398 4562 11450
rect 4624 11398 4636 11450
rect 4698 11398 4700 11450
rect 4538 11396 4562 11398
rect 4618 11396 4642 11398
rect 4698 11396 4722 11398
rect 4482 11376 4778 11396
rect 4816 11218 4844 12702
rect 5736 12306 5764 14167
rect 6840 14090 6868 14167
rect 6840 14062 7052 14090
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4482 10364 4778 10384
rect 4538 10362 4562 10364
rect 4618 10362 4642 10364
rect 4698 10362 4722 10364
rect 4560 10310 4562 10362
rect 4624 10310 4636 10362
rect 4698 10310 4700 10362
rect 4538 10308 4562 10310
rect 4618 10308 4642 10310
rect 4698 10308 4722 10310
rect 4482 10288 4778 10308
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 2719 9820 3015 9840
rect 2775 9818 2799 9820
rect 2855 9818 2879 9820
rect 2935 9818 2959 9820
rect 2797 9766 2799 9818
rect 2861 9766 2873 9818
rect 2935 9766 2937 9818
rect 2775 9764 2799 9766
rect 2855 9764 2879 9766
rect 2935 9764 2959 9766
rect 2719 9744 3015 9764
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2516 8022 2544 9114
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2719 8732 3015 8752
rect 2775 8730 2799 8732
rect 2855 8730 2879 8732
rect 2935 8730 2959 8732
rect 2797 8678 2799 8730
rect 2861 8678 2873 8730
rect 2935 8678 2937 8730
rect 2775 8676 2799 8678
rect 2855 8676 2879 8678
rect 2935 8676 2959 8678
rect 2719 8656 3015 8676
rect 2872 8492 2924 8498
rect 2700 8452 2872 8480
rect 2700 8294 2728 8452
rect 2872 8434 2924 8440
rect 3068 8430 3096 8978
rect 3436 8634 3464 9930
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3712 9042 3740 9658
rect 4080 9518 4108 10134
rect 4908 10130 4936 10474
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 8090 2820 8230
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2504 8016 2556 8022
rect 2884 7970 2912 8298
rect 2504 7958 2556 7964
rect 2700 7942 2912 7970
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 2700 7886 2728 7942
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 6225 2452 7686
rect 2719 7644 3015 7664
rect 2775 7642 2799 7644
rect 2855 7642 2879 7644
rect 2935 7642 2959 7644
rect 2797 7590 2799 7642
rect 2861 7590 2873 7642
rect 2935 7590 2937 7642
rect 2775 7588 2799 7590
rect 2855 7588 2879 7590
rect 2935 7588 2959 7590
rect 2719 7568 3015 7588
rect 2719 6556 3015 6576
rect 2775 6554 2799 6556
rect 2855 6554 2879 6556
rect 2935 6554 2959 6556
rect 2797 6502 2799 6554
rect 2861 6502 2873 6554
rect 2935 6502 2937 6554
rect 2775 6500 2799 6502
rect 2855 6500 2879 6502
rect 2935 6500 2959 6502
rect 2719 6480 3015 6500
rect 2410 6216 2466 6225
rect 2410 6151 2412 6160
rect 2464 6151 2466 6160
rect 2412 6122 2464 6128
rect 2424 6091 2452 6122
rect 3160 5778 3188 7958
rect 3252 6254 3280 8570
rect 3620 8430 3648 8774
rect 4172 8566 4200 9318
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4356 8430 4384 10066
rect 4816 9994 4844 10066
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4482 9276 4778 9296
rect 4538 9274 4562 9276
rect 4618 9274 4642 9276
rect 4698 9274 4722 9276
rect 4560 9222 4562 9274
rect 4624 9222 4636 9274
rect 4698 9222 4700 9274
rect 4538 9220 4562 9222
rect 4618 9220 4642 9222
rect 4698 9220 4722 9222
rect 4482 9200 4778 9220
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4448 8498 4476 8978
rect 5000 8634 5028 9454
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 5092 8430 5120 10202
rect 5170 10160 5226 10169
rect 5170 10095 5226 10104
rect 5184 9110 5212 10095
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5276 9722 5304 9998
rect 5460 9897 5488 12038
rect 6246 11996 6542 12016
rect 6302 11994 6326 11996
rect 6382 11994 6406 11996
rect 6462 11994 6486 11996
rect 6324 11942 6326 11994
rect 6388 11942 6400 11994
rect 6462 11942 6464 11994
rect 6302 11940 6326 11942
rect 6382 11940 6406 11942
rect 6462 11940 6486 11942
rect 6246 11920 6542 11940
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5446 9888 5502 9897
rect 5446 9823 5502 9832
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5460 9518 5488 9658
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5446 9344 5502 9353
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5276 8430 5304 9046
rect 5368 8430 5396 9318
rect 5446 9279 5502 9288
rect 5460 9042 5488 9279
rect 5552 9058 5580 11086
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 10198 5672 10610
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9518 5672 9930
rect 5632 9512 5684 9518
rect 5736 9489 5764 11494
rect 6012 10742 6040 11494
rect 7024 11286 7052 14062
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11694 7696 12038
rect 7944 11762 7972 14167
rect 8009 12540 8305 12560
rect 8065 12538 8089 12540
rect 8145 12538 8169 12540
rect 8225 12538 8249 12540
rect 8087 12486 8089 12538
rect 8151 12486 8163 12538
rect 8225 12486 8227 12538
rect 8065 12484 8089 12486
rect 8145 12484 8169 12486
rect 8225 12484 8249 12486
rect 8009 12464 8305 12484
rect 8956 12306 8984 14167
rect 10060 14090 10088 14167
rect 9692 14062 10088 14090
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7668 11218 7696 11630
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 10266 5856 10542
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 9874 5856 10066
rect 5828 9846 5948 9874
rect 5816 9512 5868 9518
rect 5632 9454 5684 9460
rect 5722 9480 5778 9489
rect 5816 9454 5868 9460
rect 5722 9415 5778 9424
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5448 9036 5500 9042
rect 5552 9030 5672 9058
rect 5448 8978 5500 8984
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 2719 5468 3015 5488
rect 2775 5466 2799 5468
rect 2855 5466 2879 5468
rect 2935 5466 2959 5468
rect 2797 5414 2799 5466
rect 2861 5414 2873 5466
rect 2935 5414 2937 5466
rect 2775 5412 2799 5414
rect 2855 5412 2879 5414
rect 2935 5412 2959 5414
rect 2719 5392 3015 5412
rect 2719 4380 3015 4400
rect 2775 4378 2799 4380
rect 2855 4378 2879 4380
rect 2935 4378 2959 4380
rect 2797 4326 2799 4378
rect 2861 4326 2873 4378
rect 2935 4326 2937 4378
rect 2775 4324 2799 4326
rect 2855 4324 2879 4326
rect 2935 4324 2959 4326
rect 2719 4304 3015 4324
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2608 800 2636 3674
rect 2719 3292 3015 3312
rect 2775 3290 2799 3292
rect 2855 3290 2879 3292
rect 2935 3290 2959 3292
rect 2797 3238 2799 3290
rect 2861 3238 2873 3290
rect 2935 3238 2937 3290
rect 2775 3236 2799 3238
rect 2855 3236 2879 3238
rect 2935 3236 2959 3238
rect 2719 3216 3015 3236
rect 2719 2204 3015 2224
rect 2775 2202 2799 2204
rect 2855 2202 2879 2204
rect 2935 2202 2959 2204
rect 2797 2150 2799 2202
rect 2861 2150 2873 2202
rect 2935 2150 2937 2202
rect 2775 2148 2799 2150
rect 2855 2148 2879 2150
rect 2935 2148 2959 2150
rect 2719 2128 3015 2148
rect 3160 1329 3188 5714
rect 3252 3777 3280 6190
rect 3238 3768 3294 3777
rect 3238 3703 3294 3712
rect 3146 1320 3202 1329
rect 3146 1255 3202 1264
rect 3620 800 3648 8026
rect 3712 7750 3740 8366
rect 5460 8294 5488 8978
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 4482 8188 4778 8208
rect 4538 8186 4562 8188
rect 4618 8186 4642 8188
rect 4698 8186 4722 8188
rect 4560 8134 4562 8186
rect 4624 8134 4636 8186
rect 4698 8134 4700 8186
rect 4538 8132 4562 8134
rect 4618 8132 4642 8134
rect 4698 8132 4722 8134
rect 4482 8112 4778 8132
rect 4436 7880 4488 7886
rect 4434 7848 4436 7857
rect 4488 7848 4490 7857
rect 4434 7783 4490 7792
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 5644 7478 5672 9030
rect 5736 8956 5764 9318
rect 5828 9178 5856 9454
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5816 8968 5868 8974
rect 5736 8928 5816 8956
rect 5816 8910 5868 8916
rect 5920 8412 5948 9846
rect 5998 9752 6054 9761
rect 5998 9687 6054 9696
rect 6012 8514 6040 9687
rect 6104 9586 6132 11154
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6246 10908 6542 10928
rect 6302 10906 6326 10908
rect 6382 10906 6406 10908
rect 6462 10906 6486 10908
rect 6324 10854 6326 10906
rect 6388 10854 6400 10906
rect 6462 10854 6464 10906
rect 6302 10852 6326 10854
rect 6382 10852 6406 10854
rect 6462 10852 6486 10854
rect 6246 10832 6542 10852
rect 6840 10606 6868 10950
rect 7668 10810 7696 11154
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6656 9874 6684 10542
rect 6840 10470 6868 10542
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6736 10124 6788 10130
rect 6840 10112 6868 10406
rect 6788 10084 6868 10112
rect 6736 10066 6788 10072
rect 6656 9846 6868 9874
rect 6246 9820 6542 9840
rect 6302 9818 6326 9820
rect 6382 9818 6406 9820
rect 6462 9818 6486 9820
rect 6324 9766 6326 9818
rect 6388 9766 6400 9818
rect 6462 9766 6464 9818
rect 6302 9764 6326 9766
rect 6382 9764 6406 9766
rect 6462 9764 6486 9766
rect 6246 9744 6542 9764
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6196 8974 6224 9114
rect 6288 9042 6316 9318
rect 6840 9178 6868 9846
rect 6932 9518 6960 10474
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7024 9042 7052 9998
rect 7300 9722 7328 10542
rect 7472 10192 7524 10198
rect 7470 10160 7472 10169
rect 7524 10160 7526 10169
rect 7470 10095 7526 10104
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7378 10024 7434 10033
rect 7378 9959 7434 9968
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 9178 7328 9454
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6184 8968 6236 8974
rect 6104 8928 6184 8956
rect 6104 8616 6132 8928
rect 6368 8968 6420 8974
rect 6184 8910 6236 8916
rect 6366 8936 6368 8945
rect 6736 8968 6788 8974
rect 6420 8936 6422 8945
rect 6736 8910 6788 8916
rect 6366 8871 6422 8880
rect 6246 8732 6542 8752
rect 6302 8730 6326 8732
rect 6382 8730 6406 8732
rect 6462 8730 6486 8732
rect 6324 8678 6326 8730
rect 6388 8678 6400 8730
rect 6462 8678 6464 8730
rect 6302 8676 6326 8678
rect 6382 8676 6406 8678
rect 6462 8676 6486 8678
rect 6246 8656 6542 8676
rect 6104 8588 6224 8616
rect 6012 8486 6132 8514
rect 6000 8424 6052 8430
rect 5920 8384 6000 8412
rect 6000 8366 6052 8372
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 4712 7336 4764 7342
rect 4896 7336 4948 7342
rect 4764 7296 4844 7324
rect 4712 7278 4764 7284
rect 4482 7100 4778 7120
rect 4538 7098 4562 7100
rect 4618 7098 4642 7100
rect 4698 7098 4722 7100
rect 4560 7046 4562 7098
rect 4624 7046 4636 7098
rect 4698 7046 4700 7098
rect 4538 7044 4562 7046
rect 4618 7044 4642 7046
rect 4698 7044 4722 7046
rect 4482 7024 4778 7044
rect 4816 6730 4844 7296
rect 4896 7278 4948 7284
rect 5446 7304 5502 7313
rect 4908 6866 4936 7278
rect 5446 7239 5502 7248
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6866 5028 7142
rect 5460 6934 5488 7239
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5644 6798 5672 7414
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 4482 6012 4778 6032
rect 4538 6010 4562 6012
rect 4618 6010 4642 6012
rect 4698 6010 4722 6012
rect 4560 5958 4562 6010
rect 4624 5958 4636 6010
rect 4698 5958 4700 6010
rect 4538 5956 4562 5958
rect 4618 5956 4642 5958
rect 4698 5956 4722 5958
rect 4482 5936 4778 5956
rect 4482 4924 4778 4944
rect 4538 4922 4562 4924
rect 4618 4922 4642 4924
rect 4698 4922 4722 4924
rect 4560 4870 4562 4922
rect 4624 4870 4636 4922
rect 4698 4870 4700 4922
rect 4538 4868 4562 4870
rect 4618 4868 4642 4870
rect 4698 4868 4722 4870
rect 4482 4848 4778 4868
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4482 3836 4778 3856
rect 4538 3834 4562 3836
rect 4618 3834 4642 3836
rect 4698 3834 4722 3836
rect 4560 3782 4562 3834
rect 4624 3782 4636 3834
rect 4698 3782 4700 3834
rect 4538 3780 4562 3782
rect 4618 3780 4642 3782
rect 4698 3780 4722 3782
rect 4482 3760 4778 3780
rect 4482 2748 4778 2768
rect 4538 2746 4562 2748
rect 4618 2746 4642 2748
rect 4698 2746 4722 2748
rect 4560 2694 4562 2746
rect 4624 2694 4636 2746
rect 4698 2694 4700 2746
rect 4538 2692 4562 2694
rect 4618 2692 4642 2694
rect 4698 2692 4722 2694
rect 4482 2672 4778 2692
rect 4816 2530 4844 4082
rect 5552 4026 5580 6666
rect 5644 4146 5672 6734
rect 5828 6322 5856 7890
rect 5920 7002 5948 8230
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6012 6934 6040 7822
rect 6104 7528 6132 8486
rect 6196 8090 6224 8588
rect 6748 8362 6776 8910
rect 6840 8566 6868 8978
rect 7024 8906 7052 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6246 7644 6542 7664
rect 6302 7642 6326 7644
rect 6382 7642 6406 7644
rect 6462 7642 6486 7644
rect 6324 7590 6326 7642
rect 6388 7590 6400 7642
rect 6462 7590 6464 7642
rect 6302 7588 6326 7590
rect 6382 7588 6406 7590
rect 6462 7588 6486 7590
rect 6246 7568 6542 7588
rect 6104 7500 6224 7528
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6104 6866 6132 7278
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5736 5574 5764 6190
rect 5920 5914 5948 6802
rect 6196 6730 6224 7500
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6656 6866 6684 7346
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 6254 6132 6598
rect 6246 6556 6542 6576
rect 6302 6554 6326 6556
rect 6382 6554 6406 6556
rect 6462 6554 6486 6556
rect 6324 6502 6326 6554
rect 6388 6502 6400 6554
rect 6462 6502 6464 6554
rect 6302 6500 6326 6502
rect 6382 6500 6406 6502
rect 6462 6500 6486 6502
rect 6246 6480 6542 6500
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6274 6352 6330 6361
rect 6274 6287 6330 6296
rect 6288 6254 6316 6287
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6748 6118 6776 7686
rect 6840 7478 6868 8502
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 7002 6868 7278
rect 6932 7206 6960 7958
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6748 5778 6776 6054
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 6246 5468 6542 5488
rect 6302 5466 6326 5468
rect 6382 5466 6406 5468
rect 6462 5466 6486 5468
rect 6324 5414 6326 5466
rect 6388 5414 6400 5466
rect 6462 5414 6464 5466
rect 6302 5412 6326 5414
rect 6382 5412 6406 5414
rect 6462 5412 6486 5414
rect 6246 5392 6542 5412
rect 6246 4380 6542 4400
rect 6302 4378 6326 4380
rect 6382 4378 6406 4380
rect 6462 4378 6486 4380
rect 6324 4326 6326 4378
rect 6388 4326 6400 4378
rect 6462 4326 6464 4378
rect 6302 4324 6326 4326
rect 6382 4324 6406 4326
rect 6462 4324 6486 4326
rect 6246 4304 6542 4324
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5552 3998 5764 4026
rect 4724 2502 4844 2530
rect 4724 800 4752 2502
rect 5736 800 5764 3998
rect 6840 3738 6868 6938
rect 6932 5778 6960 7142
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6246 3292 6542 3312
rect 6302 3290 6326 3292
rect 6382 3290 6406 3292
rect 6462 3290 6486 3292
rect 6324 3238 6326 3290
rect 6388 3238 6400 3290
rect 6462 3238 6464 3290
rect 6302 3236 6326 3238
rect 6382 3236 6406 3238
rect 6462 3236 6486 3238
rect 6246 3216 6542 3236
rect 7024 3058 7052 7822
rect 7116 6458 7144 7890
rect 7300 7546 7328 9114
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7208 3670 7236 7210
rect 7392 6254 7420 9959
rect 7668 9926 7696 10066
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7470 9616 7526 9625
rect 7470 9551 7526 9560
rect 7484 9518 7512 9551
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7668 9364 7696 9862
rect 7760 9586 7788 10610
rect 7852 10033 7880 10610
rect 7838 10024 7894 10033
rect 7838 9959 7894 9968
rect 7944 9926 7972 11562
rect 8009 11452 8305 11472
rect 8065 11450 8089 11452
rect 8145 11450 8169 11452
rect 8225 11450 8249 11452
rect 8087 11398 8089 11450
rect 8151 11398 8163 11450
rect 8225 11398 8227 11450
rect 8065 11396 8089 11398
rect 8145 11396 8169 11398
rect 8225 11396 8249 11398
rect 8009 11376 8305 11396
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8312 10810 8340 11018
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8404 10538 8432 11086
rect 9692 10742 9720 14062
rect 10690 13696 10746 13705
rect 10690 13631 10746 13640
rect 9772 11996 10068 12016
rect 9828 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 9850 11942 9852 11994
rect 9914 11942 9926 11994
rect 9988 11942 9990 11994
rect 9828 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 9772 11920 10068 11940
rect 10704 11354 10732 13631
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10782 11248 10838 11257
rect 10416 11212 10468 11218
rect 10782 11183 10838 11192
rect 10416 11154 10468 11160
rect 9772 10908 10068 10928
rect 9828 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 9850 10854 9852 10906
rect 9914 10854 9926 10906
rect 9988 10854 9990 10906
rect 9828 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 9772 10832 10068 10852
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8009 10364 8305 10384
rect 8065 10362 8089 10364
rect 8145 10362 8169 10364
rect 8225 10362 8249 10364
rect 8087 10310 8089 10362
rect 8151 10310 8163 10362
rect 8225 10310 8227 10362
rect 8065 10308 8089 10310
rect 8145 10308 8169 10310
rect 8225 10308 8249 10310
rect 8009 10288 8305 10308
rect 8404 10130 8432 10474
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7944 9722 7972 9862
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7668 9336 7788 9364
rect 7760 8974 7788 9336
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7484 8430 7512 8774
rect 7576 8566 7604 8774
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7576 8430 7604 8502
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7944 8412 7972 9454
rect 8009 9276 8305 9296
rect 8065 9274 8089 9276
rect 8145 9274 8169 9276
rect 8225 9274 8249 9276
rect 8087 9222 8089 9274
rect 8151 9222 8163 9274
rect 8225 9222 8227 9274
rect 8065 9220 8089 9222
rect 8145 9220 8169 9222
rect 8225 9220 8249 9222
rect 8009 9200 8305 9220
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8537 8248 8842
rect 8206 8528 8262 8537
rect 8206 8463 8208 8472
rect 8260 8463 8262 8472
rect 8208 8434 8260 8440
rect 8024 8424 8076 8430
rect 7944 8384 8024 8412
rect 7840 8288 7892 8294
rect 7668 8236 7840 8242
rect 7668 8230 7892 8236
rect 7668 8214 7880 8230
rect 7668 8022 7696 8214
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7546 7512 7890
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7576 6866 7604 6938
rect 7760 6934 7788 8026
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6254 7696 6598
rect 7852 6254 7880 8214
rect 7944 6866 7972 8384
rect 8024 8366 8076 8372
rect 8298 8392 8354 8401
rect 8298 8327 8300 8336
rect 8352 8327 8354 8336
rect 8300 8298 8352 8304
rect 8009 8188 8305 8208
rect 8065 8186 8089 8188
rect 8145 8186 8169 8188
rect 8225 8186 8249 8188
rect 8087 8134 8089 8186
rect 8151 8134 8163 8186
rect 8225 8134 8227 8186
rect 8065 8132 8089 8134
rect 8145 8132 8169 8134
rect 8225 8132 8249 8134
rect 8009 8112 8305 8132
rect 8404 7886 8432 10066
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8128 7342 8156 7482
rect 8220 7342 8248 7822
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8009 7100 8305 7120
rect 8065 7098 8089 7100
rect 8145 7098 8169 7100
rect 8225 7098 8249 7100
rect 8087 7046 8089 7098
rect 8151 7046 8163 7098
rect 8225 7046 8227 7098
rect 8065 7044 8089 7046
rect 8145 7044 8169 7046
rect 8225 7044 8249 7046
rect 8009 7024 8305 7044
rect 8404 7002 8432 7210
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7300 5642 7328 6122
rect 7668 5778 7696 6190
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5846 7788 6122
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7852 5778 7880 6054
rect 7944 5846 7972 6802
rect 8496 6780 8524 9930
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 8090 8616 9522
rect 8680 8906 8708 10202
rect 8772 9042 8800 10542
rect 8864 10130 8892 10678
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8864 8838 8892 10066
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8588 7313 8616 7890
rect 8574 7304 8630 7313
rect 8574 7239 8630 7248
rect 8576 6792 8628 6798
rect 8496 6752 8576 6780
rect 8576 6734 8628 6740
rect 8680 6662 8708 7890
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8772 6361 8800 7822
rect 8864 7342 8892 8230
rect 8956 7410 8984 9862
rect 9048 9518 9076 10474
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9034 9344 9090 9353
rect 9034 9279 9090 9288
rect 9048 9042 9076 9279
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9140 8974 9168 9862
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9178 9260 9454
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8864 6934 8892 7278
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8758 6352 8814 6361
rect 8758 6287 8814 6296
rect 8009 6012 8305 6032
rect 8065 6010 8089 6012
rect 8145 6010 8169 6012
rect 8225 6010 8249 6012
rect 8087 5958 8089 6010
rect 8151 5958 8163 6010
rect 8225 5958 8227 6010
rect 8065 5956 8089 5958
rect 8145 5956 8169 5958
rect 8225 5956 8249 5958
rect 8009 5936 8305 5956
rect 8956 5914 8984 6802
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 9048 5642 9076 8774
rect 9140 8634 9168 8910
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9324 8537 9352 8774
rect 9310 8528 9366 8537
rect 9310 8463 9366 8472
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 6118 9168 8366
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 7750 9352 8298
rect 9416 7857 9444 9998
rect 9494 9616 9550 9625
rect 9494 9551 9496 9560
rect 9548 9551 9550 9560
rect 9496 9522 9548 9528
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9353 9536 9386
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9508 8786 9536 9114
rect 9692 9042 9720 10406
rect 9772 9820 10068 9840
rect 9828 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 9850 9766 9852 9818
rect 9914 9766 9926 9818
rect 9988 9766 9990 9818
rect 9828 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 9772 9744 10068 9764
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9586 8936 9642 8945
rect 9784 8922 9812 8978
rect 9642 8894 9812 8922
rect 9586 8871 9642 8880
rect 9508 8758 9720 8786
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9402 7848 9458 7857
rect 9402 7783 9458 7792
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7342 9352 7686
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9312 6316 9364 6322
rect 9416 6304 9444 7783
rect 9600 7546 9628 8570
rect 9692 8498 9720 8758
rect 9772 8732 10068 8752
rect 9828 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 9850 8678 9852 8730
rect 9914 8678 9926 8730
rect 9988 8678 9990 8730
rect 9828 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 9772 8656 10068 8676
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7886 10088 8230
rect 9772 7880 9824 7886
rect 9692 7840 9772 7868
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9600 7342 9628 7482
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9692 6934 9720 7840
rect 9772 7822 9824 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9772 7644 10068 7664
rect 9828 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 9850 7590 9852 7642
rect 9914 7590 9926 7642
rect 9988 7590 9990 7642
rect 9828 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 9772 7568 10068 7588
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9784 6746 9812 7142
rect 9692 6718 9812 6746
rect 9692 6390 9720 6718
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 9772 6556 10068 6576
rect 9828 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 9850 6502 9852 6554
rect 9914 6502 9926 6554
rect 9988 6502 9990 6554
rect 9828 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 9772 6480 10068 6500
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9364 6276 9444 6304
rect 9312 6258 9364 6264
rect 9784 6254 9812 6326
rect 10152 6254 10180 6598
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8009 4924 8305 4944
rect 8065 4922 8089 4924
rect 8145 4922 8169 4924
rect 8225 4922 8249 4924
rect 8087 4870 8089 4922
rect 8151 4870 8163 4922
rect 8225 4870 8227 4922
rect 8065 4868 8089 4870
rect 8145 4868 8169 4870
rect 8225 4868 8249 4870
rect 8009 4848 8305 4868
rect 8009 3836 8305 3856
rect 8065 3834 8089 3836
rect 8145 3834 8169 3836
rect 8225 3834 8249 3836
rect 8087 3782 8089 3834
rect 8151 3782 8163 3834
rect 8225 3782 8227 3834
rect 8065 3780 8089 3782
rect 8145 3780 8169 3782
rect 8225 3780 8249 3782
rect 8009 3760 8305 3780
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7012 3052 7064 3058
rect 6840 3012 7012 3040
rect 6246 2204 6542 2224
rect 6302 2202 6326 2204
rect 6382 2202 6406 2204
rect 6462 2202 6486 2204
rect 6324 2150 6326 2202
rect 6388 2150 6400 2202
rect 6462 2150 6464 2202
rect 6302 2148 6326 2150
rect 6382 2148 6406 2150
rect 6462 2148 6486 2150
rect 6246 2128 6542 2148
rect 6840 800 6868 3012
rect 7012 2994 7064 3000
rect 7208 2514 7236 3606
rect 8009 2748 8305 2768
rect 8065 2746 8089 2748
rect 8145 2746 8169 2748
rect 8225 2746 8249 2748
rect 8087 2694 8089 2746
rect 8151 2694 8163 2746
rect 8225 2694 8227 2746
rect 8065 2692 8089 2694
rect 8145 2692 8169 2694
rect 8225 2692 8249 2694
rect 8009 2672 8305 2692
rect 8588 2514 8616 5578
rect 9232 3777 9260 6190
rect 9680 6112 9732 6118
rect 10244 6066 10272 9454
rect 10336 8430 10364 9658
rect 10324 8424 10376 8430
rect 10428 8401 10456 11154
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10520 9042 10548 9658
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9178 10640 9318
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10324 8366 10376 8372
rect 10414 8392 10470 8401
rect 10336 7954 10364 8366
rect 10414 8327 10470 8336
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10336 6934 10364 7754
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10336 6254 10364 6870
rect 10428 6390 10456 8327
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 9680 6054 9732 6060
rect 9692 5574 9720 6054
rect 10152 6038 10272 6066
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9772 5468 10068 5488
rect 9828 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 9850 5414 9852 5466
rect 9914 5414 9926 5466
rect 9988 5414 9990 5466
rect 9828 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 9772 5392 10068 5412
rect 9772 4380 10068 4400
rect 9828 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 9850 4326 9852 4378
rect 9914 4326 9926 4378
rect 9988 4326 9990 4378
rect 9828 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 9772 4304 10068 4324
rect 9218 3768 9274 3777
rect 9218 3703 9274 3712
rect 9772 3292 10068 3312
rect 9828 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 9850 3238 9852 3290
rect 9914 3238 9926 3290
rect 9988 3238 9990 3290
rect 9828 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 9772 3216 10068 3236
rect 10152 3126 10180 6038
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 3194 10272 3538
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10152 2650 10180 2926
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 7944 800 7972 2246
rect 8956 800 8984 2246
rect 9772 2204 10068 2224
rect 9828 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 9850 2150 9852 2202
rect 9914 2150 9926 2202
rect 9988 2150 9990 2202
rect 9828 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 9772 2128 10068 2148
rect 10152 1306 10180 2450
rect 10428 1329 10456 5646
rect 10520 3738 10548 8978
rect 10704 8430 10732 9590
rect 10796 9178 10824 11183
rect 11072 9518 11100 14167
rect 12176 9722 12204 14167
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7274 10640 7686
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10704 6458 10732 6802
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 6248 10652 6254
rect 10598 6216 10600 6225
rect 10652 6216 10654 6225
rect 10598 6151 10654 6160
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5710 10640 6054
rect 10704 5914 10732 6394
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5778 10824 9114
rect 10966 8800 11022 8809
rect 10966 8735 11022 8744
rect 10980 8090 11008 8735
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10060 1278 10180 1306
rect 10414 1320 10470 1329
rect 10060 800 10088 1278
rect 10414 1255 10470 1264
rect 11072 800 11100 2790
rect 12176 800 12204 3402
rect 478 0 534 800
rect 1490 0 1546 800
rect 2594 0 2650 800
rect 3606 0 3662 800
rect 4710 0 4766 800
rect 5722 0 5778 800
rect 6826 0 6882 800
rect 7930 0 7986 800
rect 8942 0 8998 800
rect 10046 0 10102 800
rect 11058 0 11114 800
rect 12162 0 12218 800
<< via2 >>
rect 3054 13640 3110 13696
rect 2719 11994 2775 11996
rect 2799 11994 2855 11996
rect 2879 11994 2935 11996
rect 2959 11994 3015 11996
rect 2719 11942 2745 11994
rect 2745 11942 2775 11994
rect 2799 11942 2809 11994
rect 2809 11942 2855 11994
rect 2879 11942 2925 11994
rect 2925 11942 2935 11994
rect 2959 11942 2989 11994
rect 2989 11942 3015 11994
rect 2719 11940 2775 11942
rect 2799 11940 2855 11942
rect 2879 11940 2935 11942
rect 2959 11940 3015 11942
rect 1398 11192 1454 11248
rect 1490 9968 1546 10024
rect 2719 10906 2775 10908
rect 2799 10906 2855 10908
rect 2879 10906 2935 10908
rect 2959 10906 3015 10908
rect 2719 10854 2745 10906
rect 2745 10854 2775 10906
rect 2799 10854 2809 10906
rect 2809 10854 2855 10906
rect 2879 10854 2925 10906
rect 2925 10854 2935 10906
rect 2959 10854 2989 10906
rect 2989 10854 3015 10906
rect 2719 10852 2775 10854
rect 2799 10852 2855 10854
rect 2879 10852 2935 10854
rect 2959 10852 3015 10854
rect 2226 8744 2282 8800
rect 4482 12538 4538 12540
rect 4562 12538 4618 12540
rect 4642 12538 4698 12540
rect 4722 12538 4778 12540
rect 4482 12486 4508 12538
rect 4508 12486 4538 12538
rect 4562 12486 4572 12538
rect 4572 12486 4618 12538
rect 4642 12486 4688 12538
rect 4688 12486 4698 12538
rect 4722 12486 4752 12538
rect 4752 12486 4778 12538
rect 4482 12484 4538 12486
rect 4562 12484 4618 12486
rect 4642 12484 4698 12486
rect 4722 12484 4778 12486
rect 4482 11450 4538 11452
rect 4562 11450 4618 11452
rect 4642 11450 4698 11452
rect 4722 11450 4778 11452
rect 4482 11398 4508 11450
rect 4508 11398 4538 11450
rect 4562 11398 4572 11450
rect 4572 11398 4618 11450
rect 4642 11398 4688 11450
rect 4688 11398 4698 11450
rect 4722 11398 4752 11450
rect 4752 11398 4778 11450
rect 4482 11396 4538 11398
rect 4562 11396 4618 11398
rect 4642 11396 4698 11398
rect 4722 11396 4778 11398
rect 4482 10362 4538 10364
rect 4562 10362 4618 10364
rect 4642 10362 4698 10364
rect 4722 10362 4778 10364
rect 4482 10310 4508 10362
rect 4508 10310 4538 10362
rect 4562 10310 4572 10362
rect 4572 10310 4618 10362
rect 4642 10310 4688 10362
rect 4688 10310 4698 10362
rect 4722 10310 4752 10362
rect 4752 10310 4778 10362
rect 4482 10308 4538 10310
rect 4562 10308 4618 10310
rect 4642 10308 4698 10310
rect 4722 10308 4778 10310
rect 2719 9818 2775 9820
rect 2799 9818 2855 9820
rect 2879 9818 2935 9820
rect 2959 9818 3015 9820
rect 2719 9766 2745 9818
rect 2745 9766 2775 9818
rect 2799 9766 2809 9818
rect 2809 9766 2855 9818
rect 2879 9766 2925 9818
rect 2925 9766 2935 9818
rect 2959 9766 2989 9818
rect 2989 9766 3015 9818
rect 2719 9764 2775 9766
rect 2799 9764 2855 9766
rect 2879 9764 2935 9766
rect 2959 9764 3015 9766
rect 2719 8730 2775 8732
rect 2799 8730 2855 8732
rect 2879 8730 2935 8732
rect 2959 8730 3015 8732
rect 2719 8678 2745 8730
rect 2745 8678 2775 8730
rect 2799 8678 2809 8730
rect 2809 8678 2855 8730
rect 2879 8678 2925 8730
rect 2925 8678 2935 8730
rect 2959 8678 2989 8730
rect 2989 8678 3015 8730
rect 2719 8676 2775 8678
rect 2799 8676 2855 8678
rect 2879 8676 2935 8678
rect 2959 8676 3015 8678
rect 2719 7642 2775 7644
rect 2799 7642 2855 7644
rect 2879 7642 2935 7644
rect 2959 7642 3015 7644
rect 2719 7590 2745 7642
rect 2745 7590 2775 7642
rect 2799 7590 2809 7642
rect 2809 7590 2855 7642
rect 2879 7590 2925 7642
rect 2925 7590 2935 7642
rect 2959 7590 2989 7642
rect 2989 7590 3015 7642
rect 2719 7588 2775 7590
rect 2799 7588 2855 7590
rect 2879 7588 2935 7590
rect 2959 7588 3015 7590
rect 2719 6554 2775 6556
rect 2799 6554 2855 6556
rect 2879 6554 2935 6556
rect 2959 6554 3015 6556
rect 2719 6502 2745 6554
rect 2745 6502 2775 6554
rect 2799 6502 2809 6554
rect 2809 6502 2855 6554
rect 2879 6502 2925 6554
rect 2925 6502 2935 6554
rect 2959 6502 2989 6554
rect 2989 6502 3015 6554
rect 2719 6500 2775 6502
rect 2799 6500 2855 6502
rect 2879 6500 2935 6502
rect 2959 6500 3015 6502
rect 2410 6180 2466 6216
rect 2410 6160 2412 6180
rect 2412 6160 2464 6180
rect 2464 6160 2466 6180
rect 4482 9274 4538 9276
rect 4562 9274 4618 9276
rect 4642 9274 4698 9276
rect 4722 9274 4778 9276
rect 4482 9222 4508 9274
rect 4508 9222 4538 9274
rect 4562 9222 4572 9274
rect 4572 9222 4618 9274
rect 4642 9222 4688 9274
rect 4688 9222 4698 9274
rect 4722 9222 4752 9274
rect 4752 9222 4778 9274
rect 4482 9220 4538 9222
rect 4562 9220 4618 9222
rect 4642 9220 4698 9222
rect 4722 9220 4778 9222
rect 5170 10104 5226 10160
rect 6246 11994 6302 11996
rect 6326 11994 6382 11996
rect 6406 11994 6462 11996
rect 6486 11994 6542 11996
rect 6246 11942 6272 11994
rect 6272 11942 6302 11994
rect 6326 11942 6336 11994
rect 6336 11942 6382 11994
rect 6406 11942 6452 11994
rect 6452 11942 6462 11994
rect 6486 11942 6516 11994
rect 6516 11942 6542 11994
rect 6246 11940 6302 11942
rect 6326 11940 6382 11942
rect 6406 11940 6462 11942
rect 6486 11940 6542 11942
rect 5446 9832 5502 9888
rect 5446 9288 5502 9344
rect 8009 12538 8065 12540
rect 8089 12538 8145 12540
rect 8169 12538 8225 12540
rect 8249 12538 8305 12540
rect 8009 12486 8035 12538
rect 8035 12486 8065 12538
rect 8089 12486 8099 12538
rect 8099 12486 8145 12538
rect 8169 12486 8215 12538
rect 8215 12486 8225 12538
rect 8249 12486 8279 12538
rect 8279 12486 8305 12538
rect 8009 12484 8065 12486
rect 8089 12484 8145 12486
rect 8169 12484 8225 12486
rect 8249 12484 8305 12486
rect 5722 9424 5778 9480
rect 2719 5466 2775 5468
rect 2799 5466 2855 5468
rect 2879 5466 2935 5468
rect 2959 5466 3015 5468
rect 2719 5414 2745 5466
rect 2745 5414 2775 5466
rect 2799 5414 2809 5466
rect 2809 5414 2855 5466
rect 2879 5414 2925 5466
rect 2925 5414 2935 5466
rect 2959 5414 2989 5466
rect 2989 5414 3015 5466
rect 2719 5412 2775 5414
rect 2799 5412 2855 5414
rect 2879 5412 2935 5414
rect 2959 5412 3015 5414
rect 2719 4378 2775 4380
rect 2799 4378 2855 4380
rect 2879 4378 2935 4380
rect 2959 4378 3015 4380
rect 2719 4326 2745 4378
rect 2745 4326 2775 4378
rect 2799 4326 2809 4378
rect 2809 4326 2855 4378
rect 2879 4326 2925 4378
rect 2925 4326 2935 4378
rect 2959 4326 2989 4378
rect 2989 4326 3015 4378
rect 2719 4324 2775 4326
rect 2799 4324 2855 4326
rect 2879 4324 2935 4326
rect 2959 4324 3015 4326
rect 2719 3290 2775 3292
rect 2799 3290 2855 3292
rect 2879 3290 2935 3292
rect 2959 3290 3015 3292
rect 2719 3238 2745 3290
rect 2745 3238 2775 3290
rect 2799 3238 2809 3290
rect 2809 3238 2855 3290
rect 2879 3238 2925 3290
rect 2925 3238 2935 3290
rect 2959 3238 2989 3290
rect 2989 3238 3015 3290
rect 2719 3236 2775 3238
rect 2799 3236 2855 3238
rect 2879 3236 2935 3238
rect 2959 3236 3015 3238
rect 2719 2202 2775 2204
rect 2799 2202 2855 2204
rect 2879 2202 2935 2204
rect 2959 2202 3015 2204
rect 2719 2150 2745 2202
rect 2745 2150 2775 2202
rect 2799 2150 2809 2202
rect 2809 2150 2855 2202
rect 2879 2150 2925 2202
rect 2925 2150 2935 2202
rect 2959 2150 2989 2202
rect 2989 2150 3015 2202
rect 2719 2148 2775 2150
rect 2799 2148 2855 2150
rect 2879 2148 2935 2150
rect 2959 2148 3015 2150
rect 3238 3712 3294 3768
rect 3146 1264 3202 1320
rect 4482 8186 4538 8188
rect 4562 8186 4618 8188
rect 4642 8186 4698 8188
rect 4722 8186 4778 8188
rect 4482 8134 4508 8186
rect 4508 8134 4538 8186
rect 4562 8134 4572 8186
rect 4572 8134 4618 8186
rect 4642 8134 4688 8186
rect 4688 8134 4698 8186
rect 4722 8134 4752 8186
rect 4752 8134 4778 8186
rect 4482 8132 4538 8134
rect 4562 8132 4618 8134
rect 4642 8132 4698 8134
rect 4722 8132 4778 8134
rect 4434 7828 4436 7848
rect 4436 7828 4488 7848
rect 4488 7828 4490 7848
rect 4434 7792 4490 7828
rect 5998 9696 6054 9752
rect 6246 10906 6302 10908
rect 6326 10906 6382 10908
rect 6406 10906 6462 10908
rect 6486 10906 6542 10908
rect 6246 10854 6272 10906
rect 6272 10854 6302 10906
rect 6326 10854 6336 10906
rect 6336 10854 6382 10906
rect 6406 10854 6452 10906
rect 6452 10854 6462 10906
rect 6486 10854 6516 10906
rect 6516 10854 6542 10906
rect 6246 10852 6302 10854
rect 6326 10852 6382 10854
rect 6406 10852 6462 10854
rect 6486 10852 6542 10854
rect 6246 9818 6302 9820
rect 6326 9818 6382 9820
rect 6406 9818 6462 9820
rect 6486 9818 6542 9820
rect 6246 9766 6272 9818
rect 6272 9766 6302 9818
rect 6326 9766 6336 9818
rect 6336 9766 6382 9818
rect 6406 9766 6452 9818
rect 6452 9766 6462 9818
rect 6486 9766 6516 9818
rect 6516 9766 6542 9818
rect 6246 9764 6302 9766
rect 6326 9764 6382 9766
rect 6406 9764 6462 9766
rect 6486 9764 6542 9766
rect 7470 10140 7472 10160
rect 7472 10140 7524 10160
rect 7524 10140 7526 10160
rect 7470 10104 7526 10140
rect 7378 9968 7434 10024
rect 6366 8916 6368 8936
rect 6368 8916 6420 8936
rect 6420 8916 6422 8936
rect 6366 8880 6422 8916
rect 6246 8730 6302 8732
rect 6326 8730 6382 8732
rect 6406 8730 6462 8732
rect 6486 8730 6542 8732
rect 6246 8678 6272 8730
rect 6272 8678 6302 8730
rect 6326 8678 6336 8730
rect 6336 8678 6382 8730
rect 6406 8678 6452 8730
rect 6452 8678 6462 8730
rect 6486 8678 6516 8730
rect 6516 8678 6542 8730
rect 6246 8676 6302 8678
rect 6326 8676 6382 8678
rect 6406 8676 6462 8678
rect 6486 8676 6542 8678
rect 4482 7098 4538 7100
rect 4562 7098 4618 7100
rect 4642 7098 4698 7100
rect 4722 7098 4778 7100
rect 4482 7046 4508 7098
rect 4508 7046 4538 7098
rect 4562 7046 4572 7098
rect 4572 7046 4618 7098
rect 4642 7046 4688 7098
rect 4688 7046 4698 7098
rect 4722 7046 4752 7098
rect 4752 7046 4778 7098
rect 4482 7044 4538 7046
rect 4562 7044 4618 7046
rect 4642 7044 4698 7046
rect 4722 7044 4778 7046
rect 5446 7248 5502 7304
rect 4482 6010 4538 6012
rect 4562 6010 4618 6012
rect 4642 6010 4698 6012
rect 4722 6010 4778 6012
rect 4482 5958 4508 6010
rect 4508 5958 4538 6010
rect 4562 5958 4572 6010
rect 4572 5958 4618 6010
rect 4642 5958 4688 6010
rect 4688 5958 4698 6010
rect 4722 5958 4752 6010
rect 4752 5958 4778 6010
rect 4482 5956 4538 5958
rect 4562 5956 4618 5958
rect 4642 5956 4698 5958
rect 4722 5956 4778 5958
rect 4482 4922 4538 4924
rect 4562 4922 4618 4924
rect 4642 4922 4698 4924
rect 4722 4922 4778 4924
rect 4482 4870 4508 4922
rect 4508 4870 4538 4922
rect 4562 4870 4572 4922
rect 4572 4870 4618 4922
rect 4642 4870 4688 4922
rect 4688 4870 4698 4922
rect 4722 4870 4752 4922
rect 4752 4870 4778 4922
rect 4482 4868 4538 4870
rect 4562 4868 4618 4870
rect 4642 4868 4698 4870
rect 4722 4868 4778 4870
rect 4482 3834 4538 3836
rect 4562 3834 4618 3836
rect 4642 3834 4698 3836
rect 4722 3834 4778 3836
rect 4482 3782 4508 3834
rect 4508 3782 4538 3834
rect 4562 3782 4572 3834
rect 4572 3782 4618 3834
rect 4642 3782 4688 3834
rect 4688 3782 4698 3834
rect 4722 3782 4752 3834
rect 4752 3782 4778 3834
rect 4482 3780 4538 3782
rect 4562 3780 4618 3782
rect 4642 3780 4698 3782
rect 4722 3780 4778 3782
rect 4482 2746 4538 2748
rect 4562 2746 4618 2748
rect 4642 2746 4698 2748
rect 4722 2746 4778 2748
rect 4482 2694 4508 2746
rect 4508 2694 4538 2746
rect 4562 2694 4572 2746
rect 4572 2694 4618 2746
rect 4642 2694 4688 2746
rect 4688 2694 4698 2746
rect 4722 2694 4752 2746
rect 4752 2694 4778 2746
rect 4482 2692 4538 2694
rect 4562 2692 4618 2694
rect 4642 2692 4698 2694
rect 4722 2692 4778 2694
rect 6246 7642 6302 7644
rect 6326 7642 6382 7644
rect 6406 7642 6462 7644
rect 6486 7642 6542 7644
rect 6246 7590 6272 7642
rect 6272 7590 6302 7642
rect 6326 7590 6336 7642
rect 6336 7590 6382 7642
rect 6406 7590 6452 7642
rect 6452 7590 6462 7642
rect 6486 7590 6516 7642
rect 6516 7590 6542 7642
rect 6246 7588 6302 7590
rect 6326 7588 6382 7590
rect 6406 7588 6462 7590
rect 6486 7588 6542 7590
rect 6246 6554 6302 6556
rect 6326 6554 6382 6556
rect 6406 6554 6462 6556
rect 6486 6554 6542 6556
rect 6246 6502 6272 6554
rect 6272 6502 6302 6554
rect 6326 6502 6336 6554
rect 6336 6502 6382 6554
rect 6406 6502 6452 6554
rect 6452 6502 6462 6554
rect 6486 6502 6516 6554
rect 6516 6502 6542 6554
rect 6246 6500 6302 6502
rect 6326 6500 6382 6502
rect 6406 6500 6462 6502
rect 6486 6500 6542 6502
rect 6274 6296 6330 6352
rect 6246 5466 6302 5468
rect 6326 5466 6382 5468
rect 6406 5466 6462 5468
rect 6486 5466 6542 5468
rect 6246 5414 6272 5466
rect 6272 5414 6302 5466
rect 6326 5414 6336 5466
rect 6336 5414 6382 5466
rect 6406 5414 6452 5466
rect 6452 5414 6462 5466
rect 6486 5414 6516 5466
rect 6516 5414 6542 5466
rect 6246 5412 6302 5414
rect 6326 5412 6382 5414
rect 6406 5412 6462 5414
rect 6486 5412 6542 5414
rect 6246 4378 6302 4380
rect 6326 4378 6382 4380
rect 6406 4378 6462 4380
rect 6486 4378 6542 4380
rect 6246 4326 6272 4378
rect 6272 4326 6302 4378
rect 6326 4326 6336 4378
rect 6336 4326 6382 4378
rect 6406 4326 6452 4378
rect 6452 4326 6462 4378
rect 6486 4326 6516 4378
rect 6516 4326 6542 4378
rect 6246 4324 6302 4326
rect 6326 4324 6382 4326
rect 6406 4324 6462 4326
rect 6486 4324 6542 4326
rect 6246 3290 6302 3292
rect 6326 3290 6382 3292
rect 6406 3290 6462 3292
rect 6486 3290 6542 3292
rect 6246 3238 6272 3290
rect 6272 3238 6302 3290
rect 6326 3238 6336 3290
rect 6336 3238 6382 3290
rect 6406 3238 6452 3290
rect 6452 3238 6462 3290
rect 6486 3238 6516 3290
rect 6516 3238 6542 3290
rect 6246 3236 6302 3238
rect 6326 3236 6382 3238
rect 6406 3236 6462 3238
rect 6486 3236 6542 3238
rect 7470 9560 7526 9616
rect 7838 9968 7894 10024
rect 8009 11450 8065 11452
rect 8089 11450 8145 11452
rect 8169 11450 8225 11452
rect 8249 11450 8305 11452
rect 8009 11398 8035 11450
rect 8035 11398 8065 11450
rect 8089 11398 8099 11450
rect 8099 11398 8145 11450
rect 8169 11398 8215 11450
rect 8215 11398 8225 11450
rect 8249 11398 8279 11450
rect 8279 11398 8305 11450
rect 8009 11396 8065 11398
rect 8089 11396 8145 11398
rect 8169 11396 8225 11398
rect 8249 11396 8305 11398
rect 10690 13640 10746 13696
rect 9772 11994 9828 11996
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 9772 11942 9798 11994
rect 9798 11942 9828 11994
rect 9852 11942 9862 11994
rect 9862 11942 9908 11994
rect 9932 11942 9978 11994
rect 9978 11942 9988 11994
rect 10012 11942 10042 11994
rect 10042 11942 10068 11994
rect 9772 11940 9828 11942
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10782 11192 10838 11248
rect 9772 10906 9828 10908
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 9772 10854 9798 10906
rect 9798 10854 9828 10906
rect 9852 10854 9862 10906
rect 9862 10854 9908 10906
rect 9932 10854 9978 10906
rect 9978 10854 9988 10906
rect 10012 10854 10042 10906
rect 10042 10854 10068 10906
rect 9772 10852 9828 10854
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 8009 10362 8065 10364
rect 8089 10362 8145 10364
rect 8169 10362 8225 10364
rect 8249 10362 8305 10364
rect 8009 10310 8035 10362
rect 8035 10310 8065 10362
rect 8089 10310 8099 10362
rect 8099 10310 8145 10362
rect 8169 10310 8215 10362
rect 8215 10310 8225 10362
rect 8249 10310 8279 10362
rect 8279 10310 8305 10362
rect 8009 10308 8065 10310
rect 8089 10308 8145 10310
rect 8169 10308 8225 10310
rect 8249 10308 8305 10310
rect 8009 9274 8065 9276
rect 8089 9274 8145 9276
rect 8169 9274 8225 9276
rect 8249 9274 8305 9276
rect 8009 9222 8035 9274
rect 8035 9222 8065 9274
rect 8089 9222 8099 9274
rect 8099 9222 8145 9274
rect 8169 9222 8215 9274
rect 8215 9222 8225 9274
rect 8249 9222 8279 9274
rect 8279 9222 8305 9274
rect 8009 9220 8065 9222
rect 8089 9220 8145 9222
rect 8169 9220 8225 9222
rect 8249 9220 8305 9222
rect 8206 8492 8262 8528
rect 8206 8472 8208 8492
rect 8208 8472 8260 8492
rect 8260 8472 8262 8492
rect 8298 8356 8354 8392
rect 8298 8336 8300 8356
rect 8300 8336 8352 8356
rect 8352 8336 8354 8356
rect 8009 8186 8065 8188
rect 8089 8186 8145 8188
rect 8169 8186 8225 8188
rect 8249 8186 8305 8188
rect 8009 8134 8035 8186
rect 8035 8134 8065 8186
rect 8089 8134 8099 8186
rect 8099 8134 8145 8186
rect 8169 8134 8215 8186
rect 8215 8134 8225 8186
rect 8249 8134 8279 8186
rect 8279 8134 8305 8186
rect 8009 8132 8065 8134
rect 8089 8132 8145 8134
rect 8169 8132 8225 8134
rect 8249 8132 8305 8134
rect 8009 7098 8065 7100
rect 8089 7098 8145 7100
rect 8169 7098 8225 7100
rect 8249 7098 8305 7100
rect 8009 7046 8035 7098
rect 8035 7046 8065 7098
rect 8089 7046 8099 7098
rect 8099 7046 8145 7098
rect 8169 7046 8215 7098
rect 8215 7046 8225 7098
rect 8249 7046 8279 7098
rect 8279 7046 8305 7098
rect 8009 7044 8065 7046
rect 8089 7044 8145 7046
rect 8169 7044 8225 7046
rect 8249 7044 8305 7046
rect 8574 7248 8630 7304
rect 9034 9288 9090 9344
rect 8758 6296 8814 6352
rect 8009 6010 8065 6012
rect 8089 6010 8145 6012
rect 8169 6010 8225 6012
rect 8249 6010 8305 6012
rect 8009 5958 8035 6010
rect 8035 5958 8065 6010
rect 8089 5958 8099 6010
rect 8099 5958 8145 6010
rect 8169 5958 8215 6010
rect 8215 5958 8225 6010
rect 8249 5958 8279 6010
rect 8279 5958 8305 6010
rect 8009 5956 8065 5958
rect 8089 5956 8145 5958
rect 8169 5956 8225 5958
rect 8249 5956 8305 5958
rect 9310 8472 9366 8528
rect 9494 9580 9550 9616
rect 9494 9560 9496 9580
rect 9496 9560 9548 9580
rect 9548 9560 9550 9580
rect 9494 9288 9550 9344
rect 9772 9818 9828 9820
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 9772 9766 9798 9818
rect 9798 9766 9828 9818
rect 9852 9766 9862 9818
rect 9862 9766 9908 9818
rect 9932 9766 9978 9818
rect 9978 9766 9988 9818
rect 10012 9766 10042 9818
rect 10042 9766 10068 9818
rect 9772 9764 9828 9766
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 9586 8880 9642 8936
rect 9402 7792 9458 7848
rect 9772 8730 9828 8732
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 9772 8678 9798 8730
rect 9798 8678 9828 8730
rect 9852 8678 9862 8730
rect 9862 8678 9908 8730
rect 9932 8678 9978 8730
rect 9978 8678 9988 8730
rect 10012 8678 10042 8730
rect 10042 8678 10068 8730
rect 9772 8676 9828 8678
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 9772 7642 9828 7644
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 9772 7590 9798 7642
rect 9798 7590 9828 7642
rect 9852 7590 9862 7642
rect 9862 7590 9908 7642
rect 9932 7590 9978 7642
rect 9978 7590 9988 7642
rect 10012 7590 10042 7642
rect 10042 7590 10068 7642
rect 9772 7588 9828 7590
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 9772 6554 9828 6556
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 9772 6502 9798 6554
rect 9798 6502 9828 6554
rect 9852 6502 9862 6554
rect 9862 6502 9908 6554
rect 9932 6502 9978 6554
rect 9978 6502 9988 6554
rect 10012 6502 10042 6554
rect 10042 6502 10068 6554
rect 9772 6500 9828 6502
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 8009 4922 8065 4924
rect 8089 4922 8145 4924
rect 8169 4922 8225 4924
rect 8249 4922 8305 4924
rect 8009 4870 8035 4922
rect 8035 4870 8065 4922
rect 8089 4870 8099 4922
rect 8099 4870 8145 4922
rect 8169 4870 8215 4922
rect 8215 4870 8225 4922
rect 8249 4870 8279 4922
rect 8279 4870 8305 4922
rect 8009 4868 8065 4870
rect 8089 4868 8145 4870
rect 8169 4868 8225 4870
rect 8249 4868 8305 4870
rect 8009 3834 8065 3836
rect 8089 3834 8145 3836
rect 8169 3834 8225 3836
rect 8249 3834 8305 3836
rect 8009 3782 8035 3834
rect 8035 3782 8065 3834
rect 8089 3782 8099 3834
rect 8099 3782 8145 3834
rect 8169 3782 8215 3834
rect 8215 3782 8225 3834
rect 8249 3782 8279 3834
rect 8279 3782 8305 3834
rect 8009 3780 8065 3782
rect 8089 3780 8145 3782
rect 8169 3780 8225 3782
rect 8249 3780 8305 3782
rect 6246 2202 6302 2204
rect 6326 2202 6382 2204
rect 6406 2202 6462 2204
rect 6486 2202 6542 2204
rect 6246 2150 6272 2202
rect 6272 2150 6302 2202
rect 6326 2150 6336 2202
rect 6336 2150 6382 2202
rect 6406 2150 6452 2202
rect 6452 2150 6462 2202
rect 6486 2150 6516 2202
rect 6516 2150 6542 2202
rect 6246 2148 6302 2150
rect 6326 2148 6382 2150
rect 6406 2148 6462 2150
rect 6486 2148 6542 2150
rect 8009 2746 8065 2748
rect 8089 2746 8145 2748
rect 8169 2746 8225 2748
rect 8249 2746 8305 2748
rect 8009 2694 8035 2746
rect 8035 2694 8065 2746
rect 8089 2694 8099 2746
rect 8099 2694 8145 2746
rect 8169 2694 8215 2746
rect 8215 2694 8225 2746
rect 8249 2694 8279 2746
rect 8279 2694 8305 2746
rect 8009 2692 8065 2694
rect 8089 2692 8145 2694
rect 8169 2692 8225 2694
rect 8249 2692 8305 2694
rect 10414 8336 10470 8392
rect 9772 5466 9828 5468
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 9772 5414 9798 5466
rect 9798 5414 9828 5466
rect 9852 5414 9862 5466
rect 9862 5414 9908 5466
rect 9932 5414 9978 5466
rect 9978 5414 9988 5466
rect 10012 5414 10042 5466
rect 10042 5414 10068 5466
rect 9772 5412 9828 5414
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 9772 4378 9828 4380
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 9772 4326 9798 4378
rect 9798 4326 9828 4378
rect 9852 4326 9862 4378
rect 9862 4326 9908 4378
rect 9932 4326 9978 4378
rect 9978 4326 9988 4378
rect 10012 4326 10042 4378
rect 10042 4326 10068 4378
rect 9772 4324 9828 4326
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 9218 3712 9274 3768
rect 9772 3290 9828 3292
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 9772 3238 9798 3290
rect 9798 3238 9828 3290
rect 9852 3238 9862 3290
rect 9862 3238 9908 3290
rect 9932 3238 9978 3290
rect 9978 3238 9988 3290
rect 10012 3238 10042 3290
rect 10042 3238 10068 3290
rect 9772 3236 9828 3238
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 9772 2202 9828 2204
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 9772 2150 9798 2202
rect 9798 2150 9828 2202
rect 9852 2150 9862 2202
rect 9862 2150 9908 2202
rect 9932 2150 9978 2202
rect 9978 2150 9988 2202
rect 10012 2150 10042 2202
rect 10042 2150 10068 2202
rect 9772 2148 9828 2150
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10598 6196 10600 6216
rect 10600 6196 10652 6216
rect 10652 6196 10654 6216
rect 10598 6160 10654 6196
rect 10966 8744 11022 8800
rect 10414 1264 10470 1320
<< metal3 >>
rect 0 13698 800 13728
rect 3049 13698 3115 13701
rect 0 13696 3115 13698
rect 0 13640 3054 13696
rect 3110 13640 3115 13696
rect 0 13638 3115 13640
rect 0 13608 800 13638
rect 3049 13635 3115 13638
rect 10685 13698 10751 13701
rect 12023 13698 12823 13728
rect 10685 13696 12823 13698
rect 10685 13640 10690 13696
rect 10746 13640 12823 13696
rect 10685 13638 12823 13640
rect 10685 13635 10751 13638
rect 12023 13608 12823 13638
rect 4470 12544 4790 12545
rect 4470 12480 4478 12544
rect 4542 12480 4558 12544
rect 4622 12480 4638 12544
rect 4702 12480 4718 12544
rect 4782 12480 4790 12544
rect 4470 12479 4790 12480
rect 7997 12544 8317 12545
rect 7997 12480 8005 12544
rect 8069 12480 8085 12544
rect 8149 12480 8165 12544
rect 8229 12480 8245 12544
rect 8309 12480 8317 12544
rect 7997 12479 8317 12480
rect 2707 12000 3027 12001
rect 2707 11936 2715 12000
rect 2779 11936 2795 12000
rect 2859 11936 2875 12000
rect 2939 11936 2955 12000
rect 3019 11936 3027 12000
rect 2707 11935 3027 11936
rect 6234 12000 6554 12001
rect 6234 11936 6242 12000
rect 6306 11936 6322 12000
rect 6386 11936 6402 12000
rect 6466 11936 6482 12000
rect 6546 11936 6554 12000
rect 6234 11935 6554 11936
rect 9760 12000 10080 12001
rect 9760 11936 9768 12000
rect 9832 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10080 12000
rect 9760 11935 10080 11936
rect 4470 11456 4790 11457
rect 4470 11392 4478 11456
rect 4542 11392 4558 11456
rect 4622 11392 4638 11456
rect 4702 11392 4718 11456
rect 4782 11392 4790 11456
rect 4470 11391 4790 11392
rect 7997 11456 8317 11457
rect 7997 11392 8005 11456
rect 8069 11392 8085 11456
rect 8149 11392 8165 11456
rect 8229 11392 8245 11456
rect 8309 11392 8317 11456
rect 7997 11391 8317 11392
rect 0 11250 800 11280
rect 1393 11250 1459 11253
rect 0 11248 1459 11250
rect 0 11192 1398 11248
rect 1454 11192 1459 11248
rect 0 11190 1459 11192
rect 0 11160 800 11190
rect 1393 11187 1459 11190
rect 10777 11250 10843 11253
rect 12023 11250 12823 11280
rect 10777 11248 12823 11250
rect 10777 11192 10782 11248
rect 10838 11192 12823 11248
rect 10777 11190 12823 11192
rect 10777 11187 10843 11190
rect 12023 11160 12823 11190
rect 2707 10912 3027 10913
rect 2707 10848 2715 10912
rect 2779 10848 2795 10912
rect 2859 10848 2875 10912
rect 2939 10848 2955 10912
rect 3019 10848 3027 10912
rect 2707 10847 3027 10848
rect 6234 10912 6554 10913
rect 6234 10848 6242 10912
rect 6306 10848 6322 10912
rect 6386 10848 6402 10912
rect 6466 10848 6482 10912
rect 6546 10848 6554 10912
rect 6234 10847 6554 10848
rect 9760 10912 10080 10913
rect 9760 10848 9768 10912
rect 9832 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10080 10912
rect 9760 10847 10080 10848
rect 4470 10368 4790 10369
rect 4470 10304 4478 10368
rect 4542 10304 4558 10368
rect 4622 10304 4638 10368
rect 4702 10304 4718 10368
rect 4782 10304 4790 10368
rect 4470 10303 4790 10304
rect 7997 10368 8317 10369
rect 7997 10304 8005 10368
rect 8069 10304 8085 10368
rect 8149 10304 8165 10368
rect 8229 10304 8245 10368
rect 8309 10304 8317 10368
rect 7997 10303 8317 10304
rect 5165 10162 5231 10165
rect 7465 10162 7531 10165
rect 5165 10160 7531 10162
rect 5165 10104 5170 10160
rect 5226 10104 7470 10160
rect 7526 10104 7531 10160
rect 5165 10102 7531 10104
rect 5165 10099 5231 10102
rect 7465 10099 7531 10102
rect 1485 10026 1551 10029
rect 7373 10026 7439 10029
rect 7833 10026 7899 10029
rect 1485 10024 7899 10026
rect 1485 9968 1490 10024
rect 1546 9968 7378 10024
rect 7434 9968 7838 10024
rect 7894 9968 7899 10024
rect 1485 9966 7899 9968
rect 1485 9963 1551 9966
rect 7373 9963 7439 9966
rect 7833 9963 7899 9966
rect 5441 9888 5507 9893
rect 5441 9832 5446 9888
rect 5502 9832 5507 9888
rect 5441 9827 5507 9832
rect 2707 9824 3027 9825
rect 2707 9760 2715 9824
rect 2779 9760 2795 9824
rect 2859 9760 2875 9824
rect 2939 9760 2955 9824
rect 3019 9760 3027 9824
rect 2707 9759 3027 9760
rect 5444 9754 5504 9827
rect 6234 9824 6554 9825
rect 6234 9760 6242 9824
rect 6306 9760 6322 9824
rect 6386 9760 6402 9824
rect 6466 9760 6482 9824
rect 6546 9760 6554 9824
rect 6234 9759 6554 9760
rect 9760 9824 10080 9825
rect 9760 9760 9768 9824
rect 9832 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10080 9824
rect 9760 9759 10080 9760
rect 5993 9754 6059 9757
rect 5444 9752 6059 9754
rect 5444 9696 5998 9752
rect 6054 9696 6059 9752
rect 5444 9694 6059 9696
rect 5993 9691 6059 9694
rect 7465 9618 7531 9621
rect 9489 9618 9555 9621
rect 7465 9616 9555 9618
rect 7465 9560 7470 9616
rect 7526 9560 9494 9616
rect 9550 9560 9555 9616
rect 7465 9558 9555 9560
rect 7465 9555 7531 9558
rect 9489 9555 9555 9558
rect 5717 9482 5783 9485
rect 5582 9480 5783 9482
rect 5582 9424 5722 9480
rect 5778 9424 5783 9480
rect 5582 9422 5783 9424
rect 5441 9346 5507 9349
rect 5582 9346 5642 9422
rect 5717 9419 5783 9422
rect 5441 9344 5642 9346
rect 5441 9288 5446 9344
rect 5502 9288 5642 9344
rect 5441 9286 5642 9288
rect 9029 9346 9095 9349
rect 9489 9346 9555 9349
rect 9029 9344 9555 9346
rect 9029 9288 9034 9344
rect 9090 9288 9494 9344
rect 9550 9288 9555 9344
rect 9029 9286 9555 9288
rect 5441 9283 5507 9286
rect 9029 9283 9095 9286
rect 9489 9283 9555 9286
rect 4470 9280 4790 9281
rect 4470 9216 4478 9280
rect 4542 9216 4558 9280
rect 4622 9216 4638 9280
rect 4702 9216 4718 9280
rect 4782 9216 4790 9280
rect 4470 9215 4790 9216
rect 7997 9280 8317 9281
rect 7997 9216 8005 9280
rect 8069 9216 8085 9280
rect 8149 9216 8165 9280
rect 8229 9216 8245 9280
rect 8309 9216 8317 9280
rect 7997 9215 8317 9216
rect 6361 8938 6427 8941
rect 9581 8938 9647 8941
rect 6361 8936 9647 8938
rect 6361 8880 6366 8936
rect 6422 8880 9586 8936
rect 9642 8880 9647 8936
rect 6361 8878 9647 8880
rect 6361 8875 6427 8878
rect 9581 8875 9647 8878
rect 0 8802 800 8832
rect 2221 8802 2287 8805
rect 0 8800 2287 8802
rect 0 8744 2226 8800
rect 2282 8744 2287 8800
rect 0 8742 2287 8744
rect 0 8712 800 8742
rect 2221 8739 2287 8742
rect 10961 8802 11027 8805
rect 12023 8802 12823 8832
rect 10961 8800 12823 8802
rect 10961 8744 10966 8800
rect 11022 8744 12823 8800
rect 10961 8742 12823 8744
rect 10961 8739 11027 8742
rect 2707 8736 3027 8737
rect 2707 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2875 8736
rect 2939 8672 2955 8736
rect 3019 8672 3027 8736
rect 2707 8671 3027 8672
rect 6234 8736 6554 8737
rect 6234 8672 6242 8736
rect 6306 8672 6322 8736
rect 6386 8672 6402 8736
rect 6466 8672 6482 8736
rect 6546 8672 6554 8736
rect 6234 8671 6554 8672
rect 9760 8736 10080 8737
rect 9760 8672 9768 8736
rect 9832 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10080 8736
rect 12023 8712 12823 8742
rect 9760 8671 10080 8672
rect 8201 8530 8267 8533
rect 9305 8530 9371 8533
rect 8201 8528 9371 8530
rect 8201 8472 8206 8528
rect 8262 8472 9310 8528
rect 9366 8472 9371 8528
rect 8201 8470 9371 8472
rect 8201 8467 8267 8470
rect 9305 8467 9371 8470
rect 8293 8394 8359 8397
rect 10409 8394 10475 8397
rect 8293 8392 10475 8394
rect 8293 8336 8298 8392
rect 8354 8336 10414 8392
rect 10470 8336 10475 8392
rect 8293 8334 10475 8336
rect 8293 8331 8359 8334
rect 10409 8331 10475 8334
rect 4470 8192 4790 8193
rect 4470 8128 4478 8192
rect 4542 8128 4558 8192
rect 4622 8128 4638 8192
rect 4702 8128 4718 8192
rect 4782 8128 4790 8192
rect 4470 8127 4790 8128
rect 7997 8192 8317 8193
rect 7997 8128 8005 8192
rect 8069 8128 8085 8192
rect 8149 8128 8165 8192
rect 8229 8128 8245 8192
rect 8309 8128 8317 8192
rect 7997 8127 8317 8128
rect 4429 7850 4495 7853
rect 9397 7850 9463 7853
rect 4429 7848 9463 7850
rect 4429 7792 4434 7848
rect 4490 7792 9402 7848
rect 9458 7792 9463 7848
rect 4429 7790 9463 7792
rect 4429 7787 4495 7790
rect 9397 7787 9463 7790
rect 2707 7648 3027 7649
rect 2707 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2875 7648
rect 2939 7584 2955 7648
rect 3019 7584 3027 7648
rect 2707 7583 3027 7584
rect 6234 7648 6554 7649
rect 6234 7584 6242 7648
rect 6306 7584 6322 7648
rect 6386 7584 6402 7648
rect 6466 7584 6482 7648
rect 6546 7584 6554 7648
rect 6234 7583 6554 7584
rect 9760 7648 10080 7649
rect 9760 7584 9768 7648
rect 9832 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10080 7648
rect 9760 7583 10080 7584
rect 5441 7306 5507 7309
rect 8569 7306 8635 7309
rect 5441 7304 8635 7306
rect 5441 7248 5446 7304
rect 5502 7248 8574 7304
rect 8630 7248 8635 7304
rect 5441 7246 8635 7248
rect 5441 7243 5507 7246
rect 8569 7243 8635 7246
rect 4470 7104 4790 7105
rect 4470 7040 4478 7104
rect 4542 7040 4558 7104
rect 4622 7040 4638 7104
rect 4702 7040 4718 7104
rect 4782 7040 4790 7104
rect 4470 7039 4790 7040
rect 7997 7104 8317 7105
rect 7997 7040 8005 7104
rect 8069 7040 8085 7104
rect 8149 7040 8165 7104
rect 8229 7040 8245 7104
rect 8309 7040 8317 7104
rect 7997 7039 8317 7040
rect 2707 6560 3027 6561
rect 2707 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2875 6560
rect 2939 6496 2955 6560
rect 3019 6496 3027 6560
rect 2707 6495 3027 6496
rect 6234 6560 6554 6561
rect 6234 6496 6242 6560
rect 6306 6496 6322 6560
rect 6386 6496 6402 6560
rect 6466 6496 6482 6560
rect 6546 6496 6554 6560
rect 6234 6495 6554 6496
rect 9760 6560 10080 6561
rect 9760 6496 9768 6560
rect 9832 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10080 6560
rect 9760 6495 10080 6496
rect 6269 6354 6335 6357
rect 8753 6354 8819 6357
rect 6269 6352 8819 6354
rect 6269 6296 6274 6352
rect 6330 6296 8758 6352
rect 8814 6296 8819 6352
rect 6269 6294 8819 6296
rect 6269 6291 6335 6294
rect 8753 6291 8819 6294
rect 0 6218 800 6248
rect 2405 6218 2471 6221
rect 0 6216 2471 6218
rect 0 6160 2410 6216
rect 2466 6160 2471 6216
rect 0 6158 2471 6160
rect 0 6128 800 6158
rect 2405 6155 2471 6158
rect 10593 6218 10659 6221
rect 12023 6218 12823 6248
rect 10593 6216 12823 6218
rect 10593 6160 10598 6216
rect 10654 6160 12823 6216
rect 10593 6158 12823 6160
rect 10593 6155 10659 6158
rect 12023 6128 12823 6158
rect 4470 6016 4790 6017
rect 4470 5952 4478 6016
rect 4542 5952 4558 6016
rect 4622 5952 4638 6016
rect 4702 5952 4718 6016
rect 4782 5952 4790 6016
rect 4470 5951 4790 5952
rect 7997 6016 8317 6017
rect 7997 5952 8005 6016
rect 8069 5952 8085 6016
rect 8149 5952 8165 6016
rect 8229 5952 8245 6016
rect 8309 5952 8317 6016
rect 7997 5951 8317 5952
rect 2707 5472 3027 5473
rect 2707 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2875 5472
rect 2939 5408 2955 5472
rect 3019 5408 3027 5472
rect 2707 5407 3027 5408
rect 6234 5472 6554 5473
rect 6234 5408 6242 5472
rect 6306 5408 6322 5472
rect 6386 5408 6402 5472
rect 6466 5408 6482 5472
rect 6546 5408 6554 5472
rect 6234 5407 6554 5408
rect 9760 5472 10080 5473
rect 9760 5408 9768 5472
rect 9832 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10080 5472
rect 9760 5407 10080 5408
rect 4470 4928 4790 4929
rect 4470 4864 4478 4928
rect 4542 4864 4558 4928
rect 4622 4864 4638 4928
rect 4702 4864 4718 4928
rect 4782 4864 4790 4928
rect 4470 4863 4790 4864
rect 7997 4928 8317 4929
rect 7997 4864 8005 4928
rect 8069 4864 8085 4928
rect 8149 4864 8165 4928
rect 8229 4864 8245 4928
rect 8309 4864 8317 4928
rect 7997 4863 8317 4864
rect 2707 4384 3027 4385
rect 2707 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2875 4384
rect 2939 4320 2955 4384
rect 3019 4320 3027 4384
rect 2707 4319 3027 4320
rect 6234 4384 6554 4385
rect 6234 4320 6242 4384
rect 6306 4320 6322 4384
rect 6386 4320 6402 4384
rect 6466 4320 6482 4384
rect 6546 4320 6554 4384
rect 6234 4319 6554 4320
rect 9760 4384 10080 4385
rect 9760 4320 9768 4384
rect 9832 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10080 4384
rect 9760 4319 10080 4320
rect 4470 3840 4790 3841
rect 0 3770 800 3800
rect 4470 3776 4478 3840
rect 4542 3776 4558 3840
rect 4622 3776 4638 3840
rect 4702 3776 4718 3840
rect 4782 3776 4790 3840
rect 4470 3775 4790 3776
rect 7997 3840 8317 3841
rect 7997 3776 8005 3840
rect 8069 3776 8085 3840
rect 8149 3776 8165 3840
rect 8229 3776 8245 3840
rect 8309 3776 8317 3840
rect 7997 3775 8317 3776
rect 3233 3770 3299 3773
rect 0 3768 3299 3770
rect 0 3712 3238 3768
rect 3294 3712 3299 3768
rect 0 3710 3299 3712
rect 0 3680 800 3710
rect 3233 3707 3299 3710
rect 9213 3770 9279 3773
rect 12023 3770 12823 3800
rect 9213 3768 12823 3770
rect 9213 3712 9218 3768
rect 9274 3712 12823 3768
rect 9213 3710 12823 3712
rect 9213 3707 9279 3710
rect 12023 3680 12823 3710
rect 2707 3296 3027 3297
rect 2707 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2875 3296
rect 2939 3232 2955 3296
rect 3019 3232 3027 3296
rect 2707 3231 3027 3232
rect 6234 3296 6554 3297
rect 6234 3232 6242 3296
rect 6306 3232 6322 3296
rect 6386 3232 6402 3296
rect 6466 3232 6482 3296
rect 6546 3232 6554 3296
rect 6234 3231 6554 3232
rect 9760 3296 10080 3297
rect 9760 3232 9768 3296
rect 9832 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10080 3296
rect 9760 3231 10080 3232
rect 4470 2752 4790 2753
rect 4470 2688 4478 2752
rect 4542 2688 4558 2752
rect 4622 2688 4638 2752
rect 4702 2688 4718 2752
rect 4782 2688 4790 2752
rect 4470 2687 4790 2688
rect 7997 2752 8317 2753
rect 7997 2688 8005 2752
rect 8069 2688 8085 2752
rect 8149 2688 8165 2752
rect 8229 2688 8245 2752
rect 8309 2688 8317 2752
rect 7997 2687 8317 2688
rect 2707 2208 3027 2209
rect 2707 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2875 2208
rect 2939 2144 2955 2208
rect 3019 2144 3027 2208
rect 2707 2143 3027 2144
rect 6234 2208 6554 2209
rect 6234 2144 6242 2208
rect 6306 2144 6322 2208
rect 6386 2144 6402 2208
rect 6466 2144 6482 2208
rect 6546 2144 6554 2208
rect 6234 2143 6554 2144
rect 9760 2208 10080 2209
rect 9760 2144 9768 2208
rect 9832 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10080 2208
rect 9760 2143 10080 2144
rect 0 1322 800 1352
rect 3141 1322 3207 1325
rect 0 1320 3207 1322
rect 0 1264 3146 1320
rect 3202 1264 3207 1320
rect 0 1262 3207 1264
rect 0 1232 800 1262
rect 3141 1259 3207 1262
rect 10409 1322 10475 1325
rect 12023 1322 12823 1352
rect 10409 1320 12823 1322
rect 10409 1264 10414 1320
rect 10470 1264 12823 1320
rect 10409 1262 12823 1264
rect 10409 1259 10475 1262
rect 12023 1232 12823 1262
<< via3 >>
rect 4478 12540 4542 12544
rect 4478 12484 4482 12540
rect 4482 12484 4538 12540
rect 4538 12484 4542 12540
rect 4478 12480 4542 12484
rect 4558 12540 4622 12544
rect 4558 12484 4562 12540
rect 4562 12484 4618 12540
rect 4618 12484 4622 12540
rect 4558 12480 4622 12484
rect 4638 12540 4702 12544
rect 4638 12484 4642 12540
rect 4642 12484 4698 12540
rect 4698 12484 4702 12540
rect 4638 12480 4702 12484
rect 4718 12540 4782 12544
rect 4718 12484 4722 12540
rect 4722 12484 4778 12540
rect 4778 12484 4782 12540
rect 4718 12480 4782 12484
rect 8005 12540 8069 12544
rect 8005 12484 8009 12540
rect 8009 12484 8065 12540
rect 8065 12484 8069 12540
rect 8005 12480 8069 12484
rect 8085 12540 8149 12544
rect 8085 12484 8089 12540
rect 8089 12484 8145 12540
rect 8145 12484 8149 12540
rect 8085 12480 8149 12484
rect 8165 12540 8229 12544
rect 8165 12484 8169 12540
rect 8169 12484 8225 12540
rect 8225 12484 8229 12540
rect 8165 12480 8229 12484
rect 8245 12540 8309 12544
rect 8245 12484 8249 12540
rect 8249 12484 8305 12540
rect 8305 12484 8309 12540
rect 8245 12480 8309 12484
rect 2715 11996 2779 12000
rect 2715 11940 2719 11996
rect 2719 11940 2775 11996
rect 2775 11940 2779 11996
rect 2715 11936 2779 11940
rect 2795 11996 2859 12000
rect 2795 11940 2799 11996
rect 2799 11940 2855 11996
rect 2855 11940 2859 11996
rect 2795 11936 2859 11940
rect 2875 11996 2939 12000
rect 2875 11940 2879 11996
rect 2879 11940 2935 11996
rect 2935 11940 2939 11996
rect 2875 11936 2939 11940
rect 2955 11996 3019 12000
rect 2955 11940 2959 11996
rect 2959 11940 3015 11996
rect 3015 11940 3019 11996
rect 2955 11936 3019 11940
rect 6242 11996 6306 12000
rect 6242 11940 6246 11996
rect 6246 11940 6302 11996
rect 6302 11940 6306 11996
rect 6242 11936 6306 11940
rect 6322 11996 6386 12000
rect 6322 11940 6326 11996
rect 6326 11940 6382 11996
rect 6382 11940 6386 11996
rect 6322 11936 6386 11940
rect 6402 11996 6466 12000
rect 6402 11940 6406 11996
rect 6406 11940 6462 11996
rect 6462 11940 6466 11996
rect 6402 11936 6466 11940
rect 6482 11996 6546 12000
rect 6482 11940 6486 11996
rect 6486 11940 6542 11996
rect 6542 11940 6546 11996
rect 6482 11936 6546 11940
rect 9768 11996 9832 12000
rect 9768 11940 9772 11996
rect 9772 11940 9828 11996
rect 9828 11940 9832 11996
rect 9768 11936 9832 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 4478 11452 4542 11456
rect 4478 11396 4482 11452
rect 4482 11396 4538 11452
rect 4538 11396 4542 11452
rect 4478 11392 4542 11396
rect 4558 11452 4622 11456
rect 4558 11396 4562 11452
rect 4562 11396 4618 11452
rect 4618 11396 4622 11452
rect 4558 11392 4622 11396
rect 4638 11452 4702 11456
rect 4638 11396 4642 11452
rect 4642 11396 4698 11452
rect 4698 11396 4702 11452
rect 4638 11392 4702 11396
rect 4718 11452 4782 11456
rect 4718 11396 4722 11452
rect 4722 11396 4778 11452
rect 4778 11396 4782 11452
rect 4718 11392 4782 11396
rect 8005 11452 8069 11456
rect 8005 11396 8009 11452
rect 8009 11396 8065 11452
rect 8065 11396 8069 11452
rect 8005 11392 8069 11396
rect 8085 11452 8149 11456
rect 8085 11396 8089 11452
rect 8089 11396 8145 11452
rect 8145 11396 8149 11452
rect 8085 11392 8149 11396
rect 8165 11452 8229 11456
rect 8165 11396 8169 11452
rect 8169 11396 8225 11452
rect 8225 11396 8229 11452
rect 8165 11392 8229 11396
rect 8245 11452 8309 11456
rect 8245 11396 8249 11452
rect 8249 11396 8305 11452
rect 8305 11396 8309 11452
rect 8245 11392 8309 11396
rect 2715 10908 2779 10912
rect 2715 10852 2719 10908
rect 2719 10852 2775 10908
rect 2775 10852 2779 10908
rect 2715 10848 2779 10852
rect 2795 10908 2859 10912
rect 2795 10852 2799 10908
rect 2799 10852 2855 10908
rect 2855 10852 2859 10908
rect 2795 10848 2859 10852
rect 2875 10908 2939 10912
rect 2875 10852 2879 10908
rect 2879 10852 2935 10908
rect 2935 10852 2939 10908
rect 2875 10848 2939 10852
rect 2955 10908 3019 10912
rect 2955 10852 2959 10908
rect 2959 10852 3015 10908
rect 3015 10852 3019 10908
rect 2955 10848 3019 10852
rect 6242 10908 6306 10912
rect 6242 10852 6246 10908
rect 6246 10852 6302 10908
rect 6302 10852 6306 10908
rect 6242 10848 6306 10852
rect 6322 10908 6386 10912
rect 6322 10852 6326 10908
rect 6326 10852 6382 10908
rect 6382 10852 6386 10908
rect 6322 10848 6386 10852
rect 6402 10908 6466 10912
rect 6402 10852 6406 10908
rect 6406 10852 6462 10908
rect 6462 10852 6466 10908
rect 6402 10848 6466 10852
rect 6482 10908 6546 10912
rect 6482 10852 6486 10908
rect 6486 10852 6542 10908
rect 6542 10852 6546 10908
rect 6482 10848 6546 10852
rect 9768 10908 9832 10912
rect 9768 10852 9772 10908
rect 9772 10852 9828 10908
rect 9828 10852 9832 10908
rect 9768 10848 9832 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 4478 10364 4542 10368
rect 4478 10308 4482 10364
rect 4482 10308 4538 10364
rect 4538 10308 4542 10364
rect 4478 10304 4542 10308
rect 4558 10364 4622 10368
rect 4558 10308 4562 10364
rect 4562 10308 4618 10364
rect 4618 10308 4622 10364
rect 4558 10304 4622 10308
rect 4638 10364 4702 10368
rect 4638 10308 4642 10364
rect 4642 10308 4698 10364
rect 4698 10308 4702 10364
rect 4638 10304 4702 10308
rect 4718 10364 4782 10368
rect 4718 10308 4722 10364
rect 4722 10308 4778 10364
rect 4778 10308 4782 10364
rect 4718 10304 4782 10308
rect 8005 10364 8069 10368
rect 8005 10308 8009 10364
rect 8009 10308 8065 10364
rect 8065 10308 8069 10364
rect 8005 10304 8069 10308
rect 8085 10364 8149 10368
rect 8085 10308 8089 10364
rect 8089 10308 8145 10364
rect 8145 10308 8149 10364
rect 8085 10304 8149 10308
rect 8165 10364 8229 10368
rect 8165 10308 8169 10364
rect 8169 10308 8225 10364
rect 8225 10308 8229 10364
rect 8165 10304 8229 10308
rect 8245 10364 8309 10368
rect 8245 10308 8249 10364
rect 8249 10308 8305 10364
rect 8305 10308 8309 10364
rect 8245 10304 8309 10308
rect 2715 9820 2779 9824
rect 2715 9764 2719 9820
rect 2719 9764 2775 9820
rect 2775 9764 2779 9820
rect 2715 9760 2779 9764
rect 2795 9820 2859 9824
rect 2795 9764 2799 9820
rect 2799 9764 2855 9820
rect 2855 9764 2859 9820
rect 2795 9760 2859 9764
rect 2875 9820 2939 9824
rect 2875 9764 2879 9820
rect 2879 9764 2935 9820
rect 2935 9764 2939 9820
rect 2875 9760 2939 9764
rect 2955 9820 3019 9824
rect 2955 9764 2959 9820
rect 2959 9764 3015 9820
rect 3015 9764 3019 9820
rect 2955 9760 3019 9764
rect 6242 9820 6306 9824
rect 6242 9764 6246 9820
rect 6246 9764 6302 9820
rect 6302 9764 6306 9820
rect 6242 9760 6306 9764
rect 6322 9820 6386 9824
rect 6322 9764 6326 9820
rect 6326 9764 6382 9820
rect 6382 9764 6386 9820
rect 6322 9760 6386 9764
rect 6402 9820 6466 9824
rect 6402 9764 6406 9820
rect 6406 9764 6462 9820
rect 6462 9764 6466 9820
rect 6402 9760 6466 9764
rect 6482 9820 6546 9824
rect 6482 9764 6486 9820
rect 6486 9764 6542 9820
rect 6542 9764 6546 9820
rect 6482 9760 6546 9764
rect 9768 9820 9832 9824
rect 9768 9764 9772 9820
rect 9772 9764 9828 9820
rect 9828 9764 9832 9820
rect 9768 9760 9832 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 4478 9276 4542 9280
rect 4478 9220 4482 9276
rect 4482 9220 4538 9276
rect 4538 9220 4542 9276
rect 4478 9216 4542 9220
rect 4558 9276 4622 9280
rect 4558 9220 4562 9276
rect 4562 9220 4618 9276
rect 4618 9220 4622 9276
rect 4558 9216 4622 9220
rect 4638 9276 4702 9280
rect 4638 9220 4642 9276
rect 4642 9220 4698 9276
rect 4698 9220 4702 9276
rect 4638 9216 4702 9220
rect 4718 9276 4782 9280
rect 4718 9220 4722 9276
rect 4722 9220 4778 9276
rect 4778 9220 4782 9276
rect 4718 9216 4782 9220
rect 8005 9276 8069 9280
rect 8005 9220 8009 9276
rect 8009 9220 8065 9276
rect 8065 9220 8069 9276
rect 8005 9216 8069 9220
rect 8085 9276 8149 9280
rect 8085 9220 8089 9276
rect 8089 9220 8145 9276
rect 8145 9220 8149 9276
rect 8085 9216 8149 9220
rect 8165 9276 8229 9280
rect 8165 9220 8169 9276
rect 8169 9220 8225 9276
rect 8225 9220 8229 9276
rect 8165 9216 8229 9220
rect 8245 9276 8309 9280
rect 8245 9220 8249 9276
rect 8249 9220 8305 9276
rect 8305 9220 8309 9276
rect 8245 9216 8309 9220
rect 2715 8732 2779 8736
rect 2715 8676 2719 8732
rect 2719 8676 2775 8732
rect 2775 8676 2779 8732
rect 2715 8672 2779 8676
rect 2795 8732 2859 8736
rect 2795 8676 2799 8732
rect 2799 8676 2855 8732
rect 2855 8676 2859 8732
rect 2795 8672 2859 8676
rect 2875 8732 2939 8736
rect 2875 8676 2879 8732
rect 2879 8676 2935 8732
rect 2935 8676 2939 8732
rect 2875 8672 2939 8676
rect 2955 8732 3019 8736
rect 2955 8676 2959 8732
rect 2959 8676 3015 8732
rect 3015 8676 3019 8732
rect 2955 8672 3019 8676
rect 6242 8732 6306 8736
rect 6242 8676 6246 8732
rect 6246 8676 6302 8732
rect 6302 8676 6306 8732
rect 6242 8672 6306 8676
rect 6322 8732 6386 8736
rect 6322 8676 6326 8732
rect 6326 8676 6382 8732
rect 6382 8676 6386 8732
rect 6322 8672 6386 8676
rect 6402 8732 6466 8736
rect 6402 8676 6406 8732
rect 6406 8676 6462 8732
rect 6462 8676 6466 8732
rect 6402 8672 6466 8676
rect 6482 8732 6546 8736
rect 6482 8676 6486 8732
rect 6486 8676 6542 8732
rect 6542 8676 6546 8732
rect 6482 8672 6546 8676
rect 9768 8732 9832 8736
rect 9768 8676 9772 8732
rect 9772 8676 9828 8732
rect 9828 8676 9832 8732
rect 9768 8672 9832 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 4478 8188 4542 8192
rect 4478 8132 4482 8188
rect 4482 8132 4538 8188
rect 4538 8132 4542 8188
rect 4478 8128 4542 8132
rect 4558 8188 4622 8192
rect 4558 8132 4562 8188
rect 4562 8132 4618 8188
rect 4618 8132 4622 8188
rect 4558 8128 4622 8132
rect 4638 8188 4702 8192
rect 4638 8132 4642 8188
rect 4642 8132 4698 8188
rect 4698 8132 4702 8188
rect 4638 8128 4702 8132
rect 4718 8188 4782 8192
rect 4718 8132 4722 8188
rect 4722 8132 4778 8188
rect 4778 8132 4782 8188
rect 4718 8128 4782 8132
rect 8005 8188 8069 8192
rect 8005 8132 8009 8188
rect 8009 8132 8065 8188
rect 8065 8132 8069 8188
rect 8005 8128 8069 8132
rect 8085 8188 8149 8192
rect 8085 8132 8089 8188
rect 8089 8132 8145 8188
rect 8145 8132 8149 8188
rect 8085 8128 8149 8132
rect 8165 8188 8229 8192
rect 8165 8132 8169 8188
rect 8169 8132 8225 8188
rect 8225 8132 8229 8188
rect 8165 8128 8229 8132
rect 8245 8188 8309 8192
rect 8245 8132 8249 8188
rect 8249 8132 8305 8188
rect 8305 8132 8309 8188
rect 8245 8128 8309 8132
rect 2715 7644 2779 7648
rect 2715 7588 2719 7644
rect 2719 7588 2775 7644
rect 2775 7588 2779 7644
rect 2715 7584 2779 7588
rect 2795 7644 2859 7648
rect 2795 7588 2799 7644
rect 2799 7588 2855 7644
rect 2855 7588 2859 7644
rect 2795 7584 2859 7588
rect 2875 7644 2939 7648
rect 2875 7588 2879 7644
rect 2879 7588 2935 7644
rect 2935 7588 2939 7644
rect 2875 7584 2939 7588
rect 2955 7644 3019 7648
rect 2955 7588 2959 7644
rect 2959 7588 3015 7644
rect 3015 7588 3019 7644
rect 2955 7584 3019 7588
rect 6242 7644 6306 7648
rect 6242 7588 6246 7644
rect 6246 7588 6302 7644
rect 6302 7588 6306 7644
rect 6242 7584 6306 7588
rect 6322 7644 6386 7648
rect 6322 7588 6326 7644
rect 6326 7588 6382 7644
rect 6382 7588 6386 7644
rect 6322 7584 6386 7588
rect 6402 7644 6466 7648
rect 6402 7588 6406 7644
rect 6406 7588 6462 7644
rect 6462 7588 6466 7644
rect 6402 7584 6466 7588
rect 6482 7644 6546 7648
rect 6482 7588 6486 7644
rect 6486 7588 6542 7644
rect 6542 7588 6546 7644
rect 6482 7584 6546 7588
rect 9768 7644 9832 7648
rect 9768 7588 9772 7644
rect 9772 7588 9828 7644
rect 9828 7588 9832 7644
rect 9768 7584 9832 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 4478 7100 4542 7104
rect 4478 7044 4482 7100
rect 4482 7044 4538 7100
rect 4538 7044 4542 7100
rect 4478 7040 4542 7044
rect 4558 7100 4622 7104
rect 4558 7044 4562 7100
rect 4562 7044 4618 7100
rect 4618 7044 4622 7100
rect 4558 7040 4622 7044
rect 4638 7100 4702 7104
rect 4638 7044 4642 7100
rect 4642 7044 4698 7100
rect 4698 7044 4702 7100
rect 4638 7040 4702 7044
rect 4718 7100 4782 7104
rect 4718 7044 4722 7100
rect 4722 7044 4778 7100
rect 4778 7044 4782 7100
rect 4718 7040 4782 7044
rect 8005 7100 8069 7104
rect 8005 7044 8009 7100
rect 8009 7044 8065 7100
rect 8065 7044 8069 7100
rect 8005 7040 8069 7044
rect 8085 7100 8149 7104
rect 8085 7044 8089 7100
rect 8089 7044 8145 7100
rect 8145 7044 8149 7100
rect 8085 7040 8149 7044
rect 8165 7100 8229 7104
rect 8165 7044 8169 7100
rect 8169 7044 8225 7100
rect 8225 7044 8229 7100
rect 8165 7040 8229 7044
rect 8245 7100 8309 7104
rect 8245 7044 8249 7100
rect 8249 7044 8305 7100
rect 8305 7044 8309 7100
rect 8245 7040 8309 7044
rect 2715 6556 2779 6560
rect 2715 6500 2719 6556
rect 2719 6500 2775 6556
rect 2775 6500 2779 6556
rect 2715 6496 2779 6500
rect 2795 6556 2859 6560
rect 2795 6500 2799 6556
rect 2799 6500 2855 6556
rect 2855 6500 2859 6556
rect 2795 6496 2859 6500
rect 2875 6556 2939 6560
rect 2875 6500 2879 6556
rect 2879 6500 2935 6556
rect 2935 6500 2939 6556
rect 2875 6496 2939 6500
rect 2955 6556 3019 6560
rect 2955 6500 2959 6556
rect 2959 6500 3015 6556
rect 3015 6500 3019 6556
rect 2955 6496 3019 6500
rect 6242 6556 6306 6560
rect 6242 6500 6246 6556
rect 6246 6500 6302 6556
rect 6302 6500 6306 6556
rect 6242 6496 6306 6500
rect 6322 6556 6386 6560
rect 6322 6500 6326 6556
rect 6326 6500 6382 6556
rect 6382 6500 6386 6556
rect 6322 6496 6386 6500
rect 6402 6556 6466 6560
rect 6402 6500 6406 6556
rect 6406 6500 6462 6556
rect 6462 6500 6466 6556
rect 6402 6496 6466 6500
rect 6482 6556 6546 6560
rect 6482 6500 6486 6556
rect 6486 6500 6542 6556
rect 6542 6500 6546 6556
rect 6482 6496 6546 6500
rect 9768 6556 9832 6560
rect 9768 6500 9772 6556
rect 9772 6500 9828 6556
rect 9828 6500 9832 6556
rect 9768 6496 9832 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 4478 6012 4542 6016
rect 4478 5956 4482 6012
rect 4482 5956 4538 6012
rect 4538 5956 4542 6012
rect 4478 5952 4542 5956
rect 4558 6012 4622 6016
rect 4558 5956 4562 6012
rect 4562 5956 4618 6012
rect 4618 5956 4622 6012
rect 4558 5952 4622 5956
rect 4638 6012 4702 6016
rect 4638 5956 4642 6012
rect 4642 5956 4698 6012
rect 4698 5956 4702 6012
rect 4638 5952 4702 5956
rect 4718 6012 4782 6016
rect 4718 5956 4722 6012
rect 4722 5956 4778 6012
rect 4778 5956 4782 6012
rect 4718 5952 4782 5956
rect 8005 6012 8069 6016
rect 8005 5956 8009 6012
rect 8009 5956 8065 6012
rect 8065 5956 8069 6012
rect 8005 5952 8069 5956
rect 8085 6012 8149 6016
rect 8085 5956 8089 6012
rect 8089 5956 8145 6012
rect 8145 5956 8149 6012
rect 8085 5952 8149 5956
rect 8165 6012 8229 6016
rect 8165 5956 8169 6012
rect 8169 5956 8225 6012
rect 8225 5956 8229 6012
rect 8165 5952 8229 5956
rect 8245 6012 8309 6016
rect 8245 5956 8249 6012
rect 8249 5956 8305 6012
rect 8305 5956 8309 6012
rect 8245 5952 8309 5956
rect 2715 5468 2779 5472
rect 2715 5412 2719 5468
rect 2719 5412 2775 5468
rect 2775 5412 2779 5468
rect 2715 5408 2779 5412
rect 2795 5468 2859 5472
rect 2795 5412 2799 5468
rect 2799 5412 2855 5468
rect 2855 5412 2859 5468
rect 2795 5408 2859 5412
rect 2875 5468 2939 5472
rect 2875 5412 2879 5468
rect 2879 5412 2935 5468
rect 2935 5412 2939 5468
rect 2875 5408 2939 5412
rect 2955 5468 3019 5472
rect 2955 5412 2959 5468
rect 2959 5412 3015 5468
rect 3015 5412 3019 5468
rect 2955 5408 3019 5412
rect 6242 5468 6306 5472
rect 6242 5412 6246 5468
rect 6246 5412 6302 5468
rect 6302 5412 6306 5468
rect 6242 5408 6306 5412
rect 6322 5468 6386 5472
rect 6322 5412 6326 5468
rect 6326 5412 6382 5468
rect 6382 5412 6386 5468
rect 6322 5408 6386 5412
rect 6402 5468 6466 5472
rect 6402 5412 6406 5468
rect 6406 5412 6462 5468
rect 6462 5412 6466 5468
rect 6402 5408 6466 5412
rect 6482 5468 6546 5472
rect 6482 5412 6486 5468
rect 6486 5412 6542 5468
rect 6542 5412 6546 5468
rect 6482 5408 6546 5412
rect 9768 5468 9832 5472
rect 9768 5412 9772 5468
rect 9772 5412 9828 5468
rect 9828 5412 9832 5468
rect 9768 5408 9832 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 4478 4924 4542 4928
rect 4478 4868 4482 4924
rect 4482 4868 4538 4924
rect 4538 4868 4542 4924
rect 4478 4864 4542 4868
rect 4558 4924 4622 4928
rect 4558 4868 4562 4924
rect 4562 4868 4618 4924
rect 4618 4868 4622 4924
rect 4558 4864 4622 4868
rect 4638 4924 4702 4928
rect 4638 4868 4642 4924
rect 4642 4868 4698 4924
rect 4698 4868 4702 4924
rect 4638 4864 4702 4868
rect 4718 4924 4782 4928
rect 4718 4868 4722 4924
rect 4722 4868 4778 4924
rect 4778 4868 4782 4924
rect 4718 4864 4782 4868
rect 8005 4924 8069 4928
rect 8005 4868 8009 4924
rect 8009 4868 8065 4924
rect 8065 4868 8069 4924
rect 8005 4864 8069 4868
rect 8085 4924 8149 4928
rect 8085 4868 8089 4924
rect 8089 4868 8145 4924
rect 8145 4868 8149 4924
rect 8085 4864 8149 4868
rect 8165 4924 8229 4928
rect 8165 4868 8169 4924
rect 8169 4868 8225 4924
rect 8225 4868 8229 4924
rect 8165 4864 8229 4868
rect 8245 4924 8309 4928
rect 8245 4868 8249 4924
rect 8249 4868 8305 4924
rect 8305 4868 8309 4924
rect 8245 4864 8309 4868
rect 2715 4380 2779 4384
rect 2715 4324 2719 4380
rect 2719 4324 2775 4380
rect 2775 4324 2779 4380
rect 2715 4320 2779 4324
rect 2795 4380 2859 4384
rect 2795 4324 2799 4380
rect 2799 4324 2855 4380
rect 2855 4324 2859 4380
rect 2795 4320 2859 4324
rect 2875 4380 2939 4384
rect 2875 4324 2879 4380
rect 2879 4324 2935 4380
rect 2935 4324 2939 4380
rect 2875 4320 2939 4324
rect 2955 4380 3019 4384
rect 2955 4324 2959 4380
rect 2959 4324 3015 4380
rect 3015 4324 3019 4380
rect 2955 4320 3019 4324
rect 6242 4380 6306 4384
rect 6242 4324 6246 4380
rect 6246 4324 6302 4380
rect 6302 4324 6306 4380
rect 6242 4320 6306 4324
rect 6322 4380 6386 4384
rect 6322 4324 6326 4380
rect 6326 4324 6382 4380
rect 6382 4324 6386 4380
rect 6322 4320 6386 4324
rect 6402 4380 6466 4384
rect 6402 4324 6406 4380
rect 6406 4324 6462 4380
rect 6462 4324 6466 4380
rect 6402 4320 6466 4324
rect 6482 4380 6546 4384
rect 6482 4324 6486 4380
rect 6486 4324 6542 4380
rect 6542 4324 6546 4380
rect 6482 4320 6546 4324
rect 9768 4380 9832 4384
rect 9768 4324 9772 4380
rect 9772 4324 9828 4380
rect 9828 4324 9832 4380
rect 9768 4320 9832 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 4478 3836 4542 3840
rect 4478 3780 4482 3836
rect 4482 3780 4538 3836
rect 4538 3780 4542 3836
rect 4478 3776 4542 3780
rect 4558 3836 4622 3840
rect 4558 3780 4562 3836
rect 4562 3780 4618 3836
rect 4618 3780 4622 3836
rect 4558 3776 4622 3780
rect 4638 3836 4702 3840
rect 4638 3780 4642 3836
rect 4642 3780 4698 3836
rect 4698 3780 4702 3836
rect 4638 3776 4702 3780
rect 4718 3836 4782 3840
rect 4718 3780 4722 3836
rect 4722 3780 4778 3836
rect 4778 3780 4782 3836
rect 4718 3776 4782 3780
rect 8005 3836 8069 3840
rect 8005 3780 8009 3836
rect 8009 3780 8065 3836
rect 8065 3780 8069 3836
rect 8005 3776 8069 3780
rect 8085 3836 8149 3840
rect 8085 3780 8089 3836
rect 8089 3780 8145 3836
rect 8145 3780 8149 3836
rect 8085 3776 8149 3780
rect 8165 3836 8229 3840
rect 8165 3780 8169 3836
rect 8169 3780 8225 3836
rect 8225 3780 8229 3836
rect 8165 3776 8229 3780
rect 8245 3836 8309 3840
rect 8245 3780 8249 3836
rect 8249 3780 8305 3836
rect 8305 3780 8309 3836
rect 8245 3776 8309 3780
rect 2715 3292 2779 3296
rect 2715 3236 2719 3292
rect 2719 3236 2775 3292
rect 2775 3236 2779 3292
rect 2715 3232 2779 3236
rect 2795 3292 2859 3296
rect 2795 3236 2799 3292
rect 2799 3236 2855 3292
rect 2855 3236 2859 3292
rect 2795 3232 2859 3236
rect 2875 3292 2939 3296
rect 2875 3236 2879 3292
rect 2879 3236 2935 3292
rect 2935 3236 2939 3292
rect 2875 3232 2939 3236
rect 2955 3292 3019 3296
rect 2955 3236 2959 3292
rect 2959 3236 3015 3292
rect 3015 3236 3019 3292
rect 2955 3232 3019 3236
rect 6242 3292 6306 3296
rect 6242 3236 6246 3292
rect 6246 3236 6302 3292
rect 6302 3236 6306 3292
rect 6242 3232 6306 3236
rect 6322 3292 6386 3296
rect 6322 3236 6326 3292
rect 6326 3236 6382 3292
rect 6382 3236 6386 3292
rect 6322 3232 6386 3236
rect 6402 3292 6466 3296
rect 6402 3236 6406 3292
rect 6406 3236 6462 3292
rect 6462 3236 6466 3292
rect 6402 3232 6466 3236
rect 6482 3292 6546 3296
rect 6482 3236 6486 3292
rect 6486 3236 6542 3292
rect 6542 3236 6546 3292
rect 6482 3232 6546 3236
rect 9768 3292 9832 3296
rect 9768 3236 9772 3292
rect 9772 3236 9828 3292
rect 9828 3236 9832 3292
rect 9768 3232 9832 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 4478 2748 4542 2752
rect 4478 2692 4482 2748
rect 4482 2692 4538 2748
rect 4538 2692 4542 2748
rect 4478 2688 4542 2692
rect 4558 2748 4622 2752
rect 4558 2692 4562 2748
rect 4562 2692 4618 2748
rect 4618 2692 4622 2748
rect 4558 2688 4622 2692
rect 4638 2748 4702 2752
rect 4638 2692 4642 2748
rect 4642 2692 4698 2748
rect 4698 2692 4702 2748
rect 4638 2688 4702 2692
rect 4718 2748 4782 2752
rect 4718 2692 4722 2748
rect 4722 2692 4778 2748
rect 4778 2692 4782 2748
rect 4718 2688 4782 2692
rect 8005 2748 8069 2752
rect 8005 2692 8009 2748
rect 8009 2692 8065 2748
rect 8065 2692 8069 2748
rect 8005 2688 8069 2692
rect 8085 2748 8149 2752
rect 8085 2692 8089 2748
rect 8089 2692 8145 2748
rect 8145 2692 8149 2748
rect 8085 2688 8149 2692
rect 8165 2748 8229 2752
rect 8165 2692 8169 2748
rect 8169 2692 8225 2748
rect 8225 2692 8229 2748
rect 8165 2688 8229 2692
rect 8245 2748 8309 2752
rect 8245 2692 8249 2748
rect 8249 2692 8305 2748
rect 8305 2692 8309 2748
rect 8245 2688 8309 2692
rect 2715 2204 2779 2208
rect 2715 2148 2719 2204
rect 2719 2148 2775 2204
rect 2775 2148 2779 2204
rect 2715 2144 2779 2148
rect 2795 2204 2859 2208
rect 2795 2148 2799 2204
rect 2799 2148 2855 2204
rect 2855 2148 2859 2204
rect 2795 2144 2859 2148
rect 2875 2204 2939 2208
rect 2875 2148 2879 2204
rect 2879 2148 2935 2204
rect 2935 2148 2939 2204
rect 2875 2144 2939 2148
rect 2955 2204 3019 2208
rect 2955 2148 2959 2204
rect 2959 2148 3015 2204
rect 3015 2148 3019 2204
rect 2955 2144 3019 2148
rect 6242 2204 6306 2208
rect 6242 2148 6246 2204
rect 6246 2148 6302 2204
rect 6302 2148 6306 2204
rect 6242 2144 6306 2148
rect 6322 2204 6386 2208
rect 6322 2148 6326 2204
rect 6326 2148 6382 2204
rect 6382 2148 6386 2204
rect 6322 2144 6386 2148
rect 6402 2204 6466 2208
rect 6402 2148 6406 2204
rect 6406 2148 6462 2204
rect 6462 2148 6466 2204
rect 6402 2144 6466 2148
rect 6482 2204 6546 2208
rect 6482 2148 6486 2204
rect 6486 2148 6542 2204
rect 6542 2148 6546 2204
rect 6482 2144 6546 2148
rect 9768 2204 9832 2208
rect 9768 2148 9772 2204
rect 9772 2148 9828 2204
rect 9828 2148 9832 2204
rect 9768 2144 9832 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
<< metal4 >>
rect 2707 12000 3027 12560
rect 2707 11936 2715 12000
rect 2779 11936 2795 12000
rect 2859 11936 2875 12000
rect 2939 11936 2955 12000
rect 3019 11936 3027 12000
rect 2707 10912 3027 11936
rect 2707 10848 2715 10912
rect 2779 10848 2795 10912
rect 2859 10848 2875 10912
rect 2939 10848 2955 10912
rect 3019 10848 3027 10912
rect 2707 9824 3027 10848
rect 2707 9760 2715 9824
rect 2779 9760 2795 9824
rect 2859 9760 2875 9824
rect 2939 9760 2955 9824
rect 3019 9760 3027 9824
rect 2707 8736 3027 9760
rect 2707 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2875 8736
rect 2939 8672 2955 8736
rect 3019 8672 3027 8736
rect 2707 7648 3027 8672
rect 2707 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2875 7648
rect 2939 7584 2955 7648
rect 3019 7584 3027 7648
rect 2707 6560 3027 7584
rect 2707 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2875 6560
rect 2939 6496 2955 6560
rect 3019 6496 3027 6560
rect 2707 5472 3027 6496
rect 2707 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2875 5472
rect 2939 5408 2955 5472
rect 3019 5408 3027 5472
rect 2707 4384 3027 5408
rect 2707 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2875 4384
rect 2939 4320 2955 4384
rect 3019 4320 3027 4384
rect 2707 3296 3027 4320
rect 2707 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2875 3296
rect 2939 3232 2955 3296
rect 3019 3232 3027 3296
rect 2707 2208 3027 3232
rect 2707 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2875 2208
rect 2939 2144 2955 2208
rect 3019 2144 3027 2208
rect 2707 2128 3027 2144
rect 4470 12544 4791 12560
rect 4470 12480 4478 12544
rect 4542 12480 4558 12544
rect 4622 12480 4638 12544
rect 4702 12480 4718 12544
rect 4782 12480 4791 12544
rect 4470 11456 4791 12480
rect 4470 11392 4478 11456
rect 4542 11392 4558 11456
rect 4622 11392 4638 11456
rect 4702 11392 4718 11456
rect 4782 11392 4791 11456
rect 4470 10368 4791 11392
rect 4470 10304 4478 10368
rect 4542 10304 4558 10368
rect 4622 10304 4638 10368
rect 4702 10304 4718 10368
rect 4782 10304 4791 10368
rect 4470 9280 4791 10304
rect 4470 9216 4478 9280
rect 4542 9216 4558 9280
rect 4622 9216 4638 9280
rect 4702 9216 4718 9280
rect 4782 9216 4791 9280
rect 4470 8192 4791 9216
rect 4470 8128 4478 8192
rect 4542 8128 4558 8192
rect 4622 8128 4638 8192
rect 4702 8128 4718 8192
rect 4782 8128 4791 8192
rect 4470 7104 4791 8128
rect 4470 7040 4478 7104
rect 4542 7040 4558 7104
rect 4622 7040 4638 7104
rect 4702 7040 4718 7104
rect 4782 7040 4791 7104
rect 4470 6016 4791 7040
rect 4470 5952 4478 6016
rect 4542 5952 4558 6016
rect 4622 5952 4638 6016
rect 4702 5952 4718 6016
rect 4782 5952 4791 6016
rect 4470 4928 4791 5952
rect 4470 4864 4478 4928
rect 4542 4864 4558 4928
rect 4622 4864 4638 4928
rect 4702 4864 4718 4928
rect 4782 4864 4791 4928
rect 4470 3840 4791 4864
rect 4470 3776 4478 3840
rect 4542 3776 4558 3840
rect 4622 3776 4638 3840
rect 4702 3776 4718 3840
rect 4782 3776 4791 3840
rect 4470 2752 4791 3776
rect 4470 2688 4478 2752
rect 4542 2688 4558 2752
rect 4622 2688 4638 2752
rect 4702 2688 4718 2752
rect 4782 2688 4791 2752
rect 4470 2128 4791 2688
rect 6234 12000 6554 12560
rect 6234 11936 6242 12000
rect 6306 11936 6322 12000
rect 6386 11936 6402 12000
rect 6466 11936 6482 12000
rect 6546 11936 6554 12000
rect 6234 10912 6554 11936
rect 6234 10848 6242 10912
rect 6306 10848 6322 10912
rect 6386 10848 6402 10912
rect 6466 10848 6482 10912
rect 6546 10848 6554 10912
rect 6234 9824 6554 10848
rect 6234 9760 6242 9824
rect 6306 9760 6322 9824
rect 6386 9760 6402 9824
rect 6466 9760 6482 9824
rect 6546 9760 6554 9824
rect 6234 8736 6554 9760
rect 6234 8672 6242 8736
rect 6306 8672 6322 8736
rect 6386 8672 6402 8736
rect 6466 8672 6482 8736
rect 6546 8672 6554 8736
rect 6234 7648 6554 8672
rect 6234 7584 6242 7648
rect 6306 7584 6322 7648
rect 6386 7584 6402 7648
rect 6466 7584 6482 7648
rect 6546 7584 6554 7648
rect 6234 6560 6554 7584
rect 6234 6496 6242 6560
rect 6306 6496 6322 6560
rect 6386 6496 6402 6560
rect 6466 6496 6482 6560
rect 6546 6496 6554 6560
rect 6234 5472 6554 6496
rect 6234 5408 6242 5472
rect 6306 5408 6322 5472
rect 6386 5408 6402 5472
rect 6466 5408 6482 5472
rect 6546 5408 6554 5472
rect 6234 4384 6554 5408
rect 6234 4320 6242 4384
rect 6306 4320 6322 4384
rect 6386 4320 6402 4384
rect 6466 4320 6482 4384
rect 6546 4320 6554 4384
rect 6234 3296 6554 4320
rect 6234 3232 6242 3296
rect 6306 3232 6322 3296
rect 6386 3232 6402 3296
rect 6466 3232 6482 3296
rect 6546 3232 6554 3296
rect 6234 2208 6554 3232
rect 6234 2144 6242 2208
rect 6306 2144 6322 2208
rect 6386 2144 6402 2208
rect 6466 2144 6482 2208
rect 6546 2144 6554 2208
rect 6234 2128 6554 2144
rect 7997 12544 8317 12560
rect 7997 12480 8005 12544
rect 8069 12480 8085 12544
rect 8149 12480 8165 12544
rect 8229 12480 8245 12544
rect 8309 12480 8317 12544
rect 7997 11456 8317 12480
rect 7997 11392 8005 11456
rect 8069 11392 8085 11456
rect 8149 11392 8165 11456
rect 8229 11392 8245 11456
rect 8309 11392 8317 11456
rect 7997 10368 8317 11392
rect 7997 10304 8005 10368
rect 8069 10304 8085 10368
rect 8149 10304 8165 10368
rect 8229 10304 8245 10368
rect 8309 10304 8317 10368
rect 7997 9280 8317 10304
rect 7997 9216 8005 9280
rect 8069 9216 8085 9280
rect 8149 9216 8165 9280
rect 8229 9216 8245 9280
rect 8309 9216 8317 9280
rect 7997 8192 8317 9216
rect 7997 8128 8005 8192
rect 8069 8128 8085 8192
rect 8149 8128 8165 8192
rect 8229 8128 8245 8192
rect 8309 8128 8317 8192
rect 7997 7104 8317 8128
rect 7997 7040 8005 7104
rect 8069 7040 8085 7104
rect 8149 7040 8165 7104
rect 8229 7040 8245 7104
rect 8309 7040 8317 7104
rect 7997 6016 8317 7040
rect 7997 5952 8005 6016
rect 8069 5952 8085 6016
rect 8149 5952 8165 6016
rect 8229 5952 8245 6016
rect 8309 5952 8317 6016
rect 7997 4928 8317 5952
rect 7997 4864 8005 4928
rect 8069 4864 8085 4928
rect 8149 4864 8165 4928
rect 8229 4864 8245 4928
rect 8309 4864 8317 4928
rect 7997 3840 8317 4864
rect 7997 3776 8005 3840
rect 8069 3776 8085 3840
rect 8149 3776 8165 3840
rect 8229 3776 8245 3840
rect 8309 3776 8317 3840
rect 7997 2752 8317 3776
rect 7997 2688 8005 2752
rect 8069 2688 8085 2752
rect 8149 2688 8165 2752
rect 8229 2688 8245 2752
rect 8309 2688 8317 2752
rect 7997 2128 8317 2688
rect 9760 12000 10081 12560
rect 9760 11936 9768 12000
rect 9832 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10081 12000
rect 9760 10912 10081 11936
rect 9760 10848 9768 10912
rect 9832 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10081 10912
rect 9760 9824 10081 10848
rect 9760 9760 9768 9824
rect 9832 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10081 9824
rect 9760 8736 10081 9760
rect 9760 8672 9768 8736
rect 9832 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10081 8736
rect 9760 7648 10081 8672
rect 9760 7584 9768 7648
rect 9832 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10081 7648
rect 9760 6560 10081 7584
rect 9760 6496 9768 6560
rect 9832 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10081 6560
rect 9760 5472 10081 6496
rect 9760 5408 9768 5472
rect 9832 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10081 5472
rect 9760 4384 10081 5408
rect 9760 4320 9768 4384
rect 9832 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10081 4384
rect 9760 3296 10081 4320
rect 9760 3232 9768 3296
rect 9832 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10081 3296
rect 9760 2208 10081 3232
rect 9760 2144 9768 2208
rect 9832 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10081 2208
rect 9760 2128 10081 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608164981
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608164981
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608164981
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608164981
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608164981
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608164981
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608164981
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608164981
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1608164981
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608164981
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1608164981
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608164981
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1608164981
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1608164981
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8188 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_82
timestamp 1608164981
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1608164981
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1608164981
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8832 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1608164981
transform 1 0 10120 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 9752 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1608164981
transform 1 0 11132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1608164981
transform 1 0 10396 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1608164981
transform 1 0 11132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101
timestamp 1608164981
transform 1 0 10396 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608164981
transform -1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608164981
transform -1 0 11684 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608164981
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608164981
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608164981
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608164981
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608164981
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1608164981
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608164981
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608164981
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608164981
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608164981
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1608164981
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1608164981
transform 1 0 11132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608164981
transform -1 0 11684 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608164981
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608164981
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608164981
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608164981
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608164981
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608164981
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608164981
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608164981
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608164981
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1608164981
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608164981
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608164981
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1608164981
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608164981
transform -1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_19
timestamp 1608164981
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_7
timestamp 1608164981
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608164981
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _150_
timestamp 1608164981
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608164981
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1608164981
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608164981
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608164981
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608164981
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608164981
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608164981
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608164981
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_111
timestamp 1608164981
transform 1 0 11316 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_105
timestamp 1608164981
transform 1 0 10764 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608164981
transform -1 0 11684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608164981
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608164981
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608164981
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608164981
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608164981
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608164981
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608164981
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608164981
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608164981
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608164981
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1608164981
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608164981
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1608164981
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608164981
transform -1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608164981
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608164981
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608164981
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608164981
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608164981
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608164981
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1608164981
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608164981
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608164981
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608164981
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608164981
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_47
timestamp 1608164981
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1608164981
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608164981
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _131_
timestamp 1608164981
transform 1 0 6072 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1608164981
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 5612 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_6_76
timestamp 1608164981
transform 1 0 8096 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608164981
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6716 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1608164981
transform 1 0 7820 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132_
timestamp 1608164981
transform 1 0 8280 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _126_
timestamp 1608164981
transform 1 0 7636 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1608164981
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1608164981
transform 1 0 8556 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1608164981
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608164981
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _121_
timestamp 1608164981
transform 1 0 9660 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _116_
timestamp 1608164981
transform 1 0 8924 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1608164981
transform 1 0 11040 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_111
timestamp 1608164981
transform 1 0 11316 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_107
timestamp 1608164981
transform 1 0 10948 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608164981
transform -1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608164981
transform -1 0 11684 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _107_
timestamp 1608164981
transform 1 0 10396 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608164981
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608164981
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608164981
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1608164981
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608164981
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608164981
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1608164981
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _130_
timestamp 1608164981
transform 1 0 5520 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 4876 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _089_
timestamp 1608164981
transform 1 0 7912 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_98
timestamp 1608164981
transform 1 0 10120 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1608164981
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608164981
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608164981
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1608164981
transform 1 0 9844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _090_
timestamp 1608164981
transform 1 0 8740 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_110
timestamp 1608164981
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608164981
transform -1 0 11684 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608164981
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608164981
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608164981
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1608164981
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_27
timestamp 1608164981
transform 1 0 3588 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1608164981
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1608164981
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _129_
timestamp 1608164981
transform 1 0 5428 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _109_
timestamp 1608164981
transform 1 0 4784 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp 1608164981
transform 1 0 7084 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608164981
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 7176 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1608164981
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1608164981
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1608164981
transform 1 0 9844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8740 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 1608164981
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1608164981
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608164981
transform -1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1608164981
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608164981
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1608164981
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1608164981
transform 1 0 2944 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608164981
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _136_
timestamp 1608164981
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  _135_
timestamp 1608164981
transform 1 0 4048 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_4  _134_
timestamp 1608164981
transform 1 0 5336 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_4  _085_
timestamp 1608164981
transform 1 0 6900 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608164981
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _133_
timestamp 1608164981
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp 1608164981
transform 1 0 11132 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608164981
transform -1 0 11684 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _149_
timestamp 1608164981
transform 1 0 10764 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1608164981
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1608164981
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608164981
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _118_
timestamp 1608164981
transform 1 0 1656 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1608164981
transform 1 0 2944 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _147_
timestamp 1608164981
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1608164981
transform 1 0 3312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _097_
timestamp 1608164981
transform 1 0 4416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 5520 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608164981
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _140_
timestamp 1608164981
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _115_
timestamp 1608164981
transform 1 0 6808 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_4  _141_
timestamp 1608164981
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1608164981
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608164981
transform -1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _080_
timestamp 1608164981
transform 1 0 10580 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_15
timestamp 1608164981
transform 1 0 2484 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1608164981
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608164981
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608164981
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _148_
timestamp 1608164981
transform 1 0 1840 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1608164981
transform 1 0 2208 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1608164981
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1608164981
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608164981
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1608164981
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _112_
timestamp 1608164981
transform 1 0 4232 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1608164981
transform 1 0 3404 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _120_
timestamp 1608164981
transform 1 0 6348 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_4  _074_
timestamp 1608164981
transform 1 0 5060 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _099_
timestamp 1608164981
transform 1 0 7912 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608164981
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608164981
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _095_
timestamp 1608164981
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608164981
transform 1 0 9016 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1608164981
transform 1 0 11040 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608164981
transform -1 0 11684 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1608164981
transform 1 0 10764 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1608164981
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp 1608164981
transform 1 0 2116 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1608164981
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_18
timestamp 1608164981
transform 1 0 2760 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_6
timestamp 1608164981
transform 1 0 1656 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608164981
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608164981
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1608164981
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _101_
timestamp 1608164981
transform 1 0 2392 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608164981
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_21
timestamp 1608164981
transform 1 0 3036 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_26
timestamp 1608164981
transform 1 0 3496 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1608164981
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1608164981
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608164981
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608164981
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1608164981
transform 1 0 4048 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1608164981
transform 1 0 4508 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _076_
timestamp 1608164981
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _145_
timestamp 1608164981
transform 1 0 4784 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _077_
timestamp 1608164981
transform 1 0 5152 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_4  _066_
timestamp 1608164981
transform 1 0 5612 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608164981
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _142_
timestamp 1608164981
transform 1 0 8096 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _123_
timestamp 1608164981
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _122_
timestamp 1608164981
transform 1 0 6808 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _071_
timestamp 1608164981
transform 1 0 6808 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1608164981
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608164981
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1608164981
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608164981
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _075_
timestamp 1608164981
transform 1 0 8740 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _072_
timestamp 1608164981
transform 1 0 9200 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1608164981
transform 1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1608164981
transform 1 0 11316 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_105
timestamp 1608164981
transform 1 0 10764 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1608164981
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608164981
transform -1 0 11684 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608164981
transform -1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608164981
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608164981
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608164981
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1608164981
transform 1 0 4692 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608164981
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1608164981
transform 1 0 5244 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _102_
timestamp 1608164981
transform 1 0 5336 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _067_
timestamp 1608164981
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608164981
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _098_
timestamp 1608164981
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _083_
timestamp 1608164981
transform 1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_92
timestamp 1608164981
transform 1 0 9568 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_80
timestamp 1608164981
transform 1 0 8464 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1608164981
transform 1 0 10672 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608164981
transform -1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608164981
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608164981
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608164981
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608164981
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608164981
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1608164981
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1608164981
transform 1 0 6164 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1608164981
transform 1 0 5796 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1608164981
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1608164981
transform 1 0 7912 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6716 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1608164981
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1608164981
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608164981
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_106
timestamp 1608164981
transform 1 0 10856 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_101
timestamp 1608164981
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608164981
transform -1 0 11684 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1608164981
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1608164981
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608164981
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608164981
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _155_
timestamp 1608164981
transform 1 0 2668 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _154_
timestamp 1608164981
transform 1 0 4416 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_17_55
timestamp 1608164981
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_77
timestamp 1608164981
transform 1 0 8188 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1608164981
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608164981
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _091_
timestamp 1608164981
transform 1 0 7544 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_89
timestamp 1608164981
transform 1 0 9292 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1608164981
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1608164981
transform 1 0 10396 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608164981
transform -1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608164981
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608164981
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608164981
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1608164981
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1608164981
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608164981
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608164981
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _152_
timestamp 1608164981
transform 1 0 4508 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_18_56
timestamp 1608164981
transform 1 0 6256 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1608164981
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_63
timestamp 1608164981
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608164981
transform 1 0 6808 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1608164981
transform 1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_94
timestamp 1608164981
transform 1 0 9752 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_92
timestamp 1608164981
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1608164981
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608164981
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_106
timestamp 1608164981
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608164981
transform -1 0 11684 0 -1 12512
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5722 14167 5778 14967 6 cbitin[0]
port 0 nsew signal input
rlabel metal2 s 4710 14167 4766 14967 6 cbitin[1]
port 1 nsew signal input
rlabel metal2 s 3606 14167 3662 14967 6 cbitin[2]
port 2 nsew signal input
rlabel metal2 s 2594 14167 2650 14967 6 cbitin[3]
port 3 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 cbitout[0]
port 4 nsew signal tristate
rlabel metal2 s 4710 0 4766 800 6 cbitout[1]
port 5 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 cbitout[2]
port 6 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 cbitout[3]
port 7 nsew signal tristate
rlabel metal2 s 1490 14167 1546 14967 6 confclk
port 8 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 confclko
port 9 nsew signal tristate
rlabel metal2 s 10046 0 10102 800 6 dempty
port 10 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 din[0]
port 11 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 din[1]
port 12 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 dout[0]
port 13 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 dout[1]
port 14 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 hempty
port 15 nsew signal tristate
rlabel metal3 s 12023 8712 12823 8832 6 hempty2
port 16 nsew signal tristate
rlabel metal3 s 0 8712 800 8832 6 lempty
port 17 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 lin[0]
port 18 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 lin[1]
port 19 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 lout[0]
port 20 nsew signal tristate
rlabel metal3 s 0 1232 800 1352 6 lout[1]
port 21 nsew signal tristate
rlabel metal3 s 12023 6128 12823 6248 6 rempty
port 22 nsew signal input
rlabel metal2 s 478 14167 534 14967 6 reset
port 23 nsew signal input
rlabel metal2 s 478 0 534 800 6 reseto
port 24 nsew signal tristate
rlabel metal3 s 12023 3680 12823 3800 6 rin[0]
port 25 nsew signal input
rlabel metal3 s 12023 1232 12823 1352 6 rin[1]
port 26 nsew signal input
rlabel metal3 s 12023 13608 12823 13728 6 rout[0]
port 27 nsew signal tristate
rlabel metal3 s 12023 11160 12823 11280 6 rout[1]
port 28 nsew signal tristate
rlabel metal2 s 8942 14167 8998 14967 6 uempty
port 29 nsew signal input
rlabel metal2 s 7930 14167 7986 14967 6 uin[0]
port 30 nsew signal input
rlabel metal2 s 6826 14167 6882 14967 6 uin[1]
port 31 nsew signal input
rlabel metal2 s 12162 14167 12218 14967 6 uout[0]
port 32 nsew signal tristate
rlabel metal2 s 11058 14167 11114 14967 6 uout[1]
port 33 nsew signal tristate
rlabel metal2 s 10046 14167 10102 14967 6 vempty
port 34 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 vempty2
port 35 nsew signal tristate
rlabel metal4 s 9761 2128 10081 12560 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 6234 2128 6554 12560 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 2707 2128 3027 12560 6 vccd1
port 38 nsew power bidirectional
rlabel metal4 s 7997 2128 8317 12560 6 vssd1
port 39 nsew ground bidirectional
rlabel metal4 s 4471 2128 4791 12560 6 vssd1
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12823 14967
<< end >>
