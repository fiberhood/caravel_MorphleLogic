magic
tech sky130A
magscale 1 2
timestamp 1608250781
<< obsli1 >>
rect 1104 2159 11684 12529
<< obsm1 >>
rect 474 2128 12222 12560
<< metal2 >>
rect 478 14167 534 14967
rect 1490 14167 1546 14967
rect 2594 14167 2650 14967
rect 3606 14167 3662 14967
rect 4710 14167 4766 14967
rect 5722 14167 5778 14967
rect 6826 14167 6882 14967
rect 7930 14167 7986 14967
rect 8942 14167 8998 14967
rect 10046 14167 10102 14967
rect 11058 14167 11114 14967
rect 12162 14167 12218 14967
rect 478 0 534 800
rect 1490 0 1546 800
rect 2594 0 2650 800
rect 3606 0 3662 800
rect 4710 0 4766 800
rect 5722 0 5778 800
rect 6826 0 6882 800
rect 7930 0 7986 800
rect 8942 0 8998 800
rect 10046 0 10102 800
rect 11058 0 11114 800
rect 12162 0 12218 800
<< obsm2 >>
rect 590 14111 1434 14167
rect 1602 14111 2538 14167
rect 2706 14111 3550 14167
rect 3718 14111 4654 14167
rect 4822 14111 5666 14167
rect 5834 14111 6770 14167
rect 6938 14111 7874 14167
rect 8042 14111 8886 14167
rect 9054 14111 9990 14167
rect 10158 14111 11002 14167
rect 11170 14111 12106 14167
rect 480 856 12216 14111
rect 590 800 1434 856
rect 1602 800 2538 856
rect 2706 800 3550 856
rect 3718 800 4654 856
rect 4822 800 5666 856
rect 5834 800 6770 856
rect 6938 800 7874 856
rect 8042 800 8886 856
rect 9054 800 9990 856
rect 10158 800 11002 856
rect 11170 800 12106 856
<< metal3 >>
rect 0 13608 800 13728
rect 12023 13608 12823 13728
rect 0 11160 800 11280
rect 12023 11160 12823 11280
rect 0 8712 800 8832
rect 12023 8712 12823 8832
rect 0 6128 800 6248
rect 12023 6128 12823 6248
rect 0 3680 800 3800
rect 12023 3680 12823 3800
rect 0 1232 800 1352
rect 12023 1232 12823 1352
<< obsm3 >>
rect 880 13528 11943 13701
rect 800 11360 12023 13528
rect 880 11080 11943 11360
rect 800 8912 12023 11080
rect 880 8632 11943 8912
rect 800 6328 12023 8632
rect 880 6048 11943 6328
rect 800 3880 12023 6048
rect 880 3600 11943 3880
rect 800 1432 12023 3600
rect 880 1259 11943 1432
<< metal4 >>
rect 2707 2128 3027 12560
rect 4471 2128 4791 12560
rect 6234 2128 6554 12560
rect 7997 2128 8317 12560
rect 9761 2128 10081 12560
<< obsm4 >>
rect 4871 2128 6154 12560
rect 6634 2128 7917 12560
rect 8397 2128 9681 12560
<< labels >>
rlabel metal2 s 5722 14167 5778 14967 6 cbitin[0]
port 1 nsew signal input
rlabel metal2 s 4710 14167 4766 14967 6 cbitin[1]
port 2 nsew signal input
rlabel metal2 s 3606 14167 3662 14967 6 cbitin[2]
port 3 nsew signal input
rlabel metal2 s 2594 14167 2650 14967 6 cbitin[3]
port 4 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 cbitout[0]
port 5 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 cbitout[1]
port 6 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 cbitout[2]
port 7 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 cbitout[3]
port 8 nsew signal output
rlabel metal2 s 1490 14167 1546 14967 6 confclk
port 9 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 confclko
port 10 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 dempty
port 11 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 din[0]
port 12 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 din[1]
port 13 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 dout[0]
port 14 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 dout[1]
port 15 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 hempty
port 16 nsew signal output
rlabel metal3 s 12023 8712 12823 8832 6 hempty2
port 17 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 lempty
port 18 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 lin[0]
port 19 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 lin[1]
port 20 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 lout[0]
port 21 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 lout[1]
port 22 nsew signal output
rlabel metal3 s 12023 6128 12823 6248 6 rempty
port 23 nsew signal input
rlabel metal2 s 478 14167 534 14967 6 reset
port 24 nsew signal input
rlabel metal2 s 478 0 534 800 6 reseto
port 25 nsew signal output
rlabel metal3 s 12023 3680 12823 3800 6 rin[0]
port 26 nsew signal input
rlabel metal3 s 12023 1232 12823 1352 6 rin[1]
port 27 nsew signal input
rlabel metal3 s 12023 13608 12823 13728 6 rout[0]
port 28 nsew signal output
rlabel metal3 s 12023 11160 12823 11280 6 rout[1]
port 29 nsew signal output
rlabel metal2 s 8942 14167 8998 14967 6 uempty
port 30 nsew signal input
rlabel metal2 s 7930 14167 7986 14967 6 uin[0]
port 31 nsew signal input
rlabel metal2 s 6826 14167 6882 14967 6 uin[1]
port 32 nsew signal input
rlabel metal2 s 12162 14167 12218 14967 6 uout[0]
port 33 nsew signal output
rlabel metal2 s 11058 14167 11114 14967 6 uout[1]
port 34 nsew signal output
rlabel metal2 s 10046 14167 10102 14967 6 vempty
port 35 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 vempty2
port 36 nsew signal output
rlabel metal4 s 9761 2128 10081 12560 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 6234 2128 6554 12560 6 vccd1
port 38 nsew power bidirectional
rlabel metal4 s 2707 2128 3027 12560 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 7997 2128 8317 12560 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 4471 2128 4791 12560 6 vssd1
port 41 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 12823 14967
string LEFview TRUE
<< end >>
